magic
tech sky130A
magscale 1 2
timestamp 1630051267
<< viali >>
rect 2513 9061 2547 9095
rect 3157 8993 3191 9027
rect 7665 8993 7699 9027
rect 1777 8925 1811 8959
rect 5733 8925 5767 8959
rect 6469 8925 6503 8959
rect 2973 8857 3007 8891
rect 5488 8857 5522 8891
rect 1961 8789 1995 8823
rect 2881 8789 2915 8823
rect 4353 8789 4387 8823
rect 6653 8789 6687 8823
rect 7113 8789 7147 8823
rect 7481 8789 7515 8823
rect 7573 8789 7607 8823
rect 2329 8585 2363 8619
rect 6377 8585 6411 8619
rect 6837 8585 6871 8619
rect 1593 8517 1627 8551
rect 1777 8517 1811 8551
rect 4712 8517 4746 8551
rect 3453 8449 3487 8483
rect 4445 8449 4479 8483
rect 6745 8449 6779 8483
rect 7849 8449 7883 8483
rect 3709 8381 3743 8415
rect 6929 8381 6963 8415
rect 5825 8313 5859 8347
rect 7665 8245 7699 8279
rect 1869 8041 1903 8075
rect 3801 8041 3835 8075
rect 6561 8041 6595 8075
rect 7665 8041 7699 8075
rect 3249 7905 3283 7939
rect 4353 7905 4387 7939
rect 2982 7837 3016 7871
rect 4169 7837 4203 7871
rect 7849 7837 7883 7871
rect 5273 7769 5307 7803
rect 4261 7701 4295 7735
rect 5365 7497 5399 7531
rect 6377 7497 6411 7531
rect 6837 7497 6871 7531
rect 2320 7429 2354 7463
rect 2053 7361 2087 7395
rect 4077 7361 4111 7395
rect 6745 7361 6779 7395
rect 6929 7293 6963 7327
rect 3433 7157 3467 7191
rect 7113 6953 7147 6987
rect 5733 6817 5767 6851
rect 3249 6749 3283 6783
rect 3893 6749 3927 6783
rect 2982 6681 3016 6715
rect 4160 6681 4194 6715
rect 6000 6681 6034 6715
rect 1869 6613 1903 6647
rect 5273 6613 5307 6647
rect 2881 6409 2915 6443
rect 3249 6409 3283 6443
rect 6377 6409 6411 6443
rect 3341 6341 3375 6375
rect 4445 6273 4479 6307
rect 4712 6273 4746 6307
rect 6745 6273 6779 6307
rect 7849 6273 7883 6307
rect 3525 6205 3559 6239
rect 6837 6205 6871 6239
rect 7021 6205 7055 6239
rect 5825 6069 5859 6103
rect 7665 6069 7699 6103
rect 5181 5865 5215 5899
rect 6377 5865 6411 5899
rect 5825 5729 5859 5763
rect 3801 5661 3835 5695
rect 6009 5661 6043 5695
rect 3249 5593 3283 5627
rect 4068 5593 4102 5627
rect 1961 5525 1995 5559
rect 5917 5525 5951 5559
rect 2053 5321 2087 5355
rect 2421 5321 2455 5355
rect 4261 5321 4295 5355
rect 5089 5321 5123 5355
rect 3126 5253 3160 5287
rect 5181 5185 5215 5219
rect 1777 5117 1811 5151
rect 1961 5117 1995 5151
rect 2881 5117 2915 5151
rect 5273 5117 5307 5151
rect 4721 5049 4755 5083
rect 4997 4777 5031 4811
rect 5181 4573 5215 4607
rect 5273 4573 5307 4607
rect 1777 4097 1811 4131
rect 1961 3961 1995 3995
rect 7665 3145 7699 3179
rect 7849 3009 7883 3043
rect 1961 2601 1995 2635
rect 2881 2601 2915 2635
rect 5641 2601 5675 2635
rect 7481 2601 7515 2635
rect 1777 2397 1811 2431
rect 2697 2397 2731 2431
rect 5457 2397 5491 2431
rect 7757 2329 7791 2363
<< metal1 >>
rect 1104 9274 8556 9296
rect 1104 9222 2224 9274
rect 2276 9222 2288 9274
rect 2340 9222 2352 9274
rect 2404 9222 2416 9274
rect 2468 9222 4708 9274
rect 4760 9222 4772 9274
rect 4824 9222 4836 9274
rect 4888 9222 4900 9274
rect 4952 9222 7192 9274
rect 7244 9222 7256 9274
rect 7308 9222 7320 9274
rect 7372 9222 7384 9274
rect 7436 9222 8556 9274
rect 1104 9200 8556 9222
rect 5534 9120 5540 9172
rect 5592 9160 5598 9172
rect 5592 9132 6500 9160
rect 5592 9120 5598 9132
rect 2501 9095 2559 9101
rect 2501 9061 2513 9095
rect 2547 9092 2559 9095
rect 2958 9092 2964 9104
rect 2547 9064 2964 9092
rect 2547 9061 2559 9064
rect 2501 9055 2559 9061
rect 2958 9052 2964 9064
rect 3016 9052 3022 9104
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 4338 9024 4344 9036
rect 3191 8996 4344 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 4338 8984 4344 8996
rect 4396 8984 4402 9036
rect 1762 8956 1768 8968
rect 1723 8928 1768 8956
rect 1762 8916 1768 8928
rect 1820 8916 1826 8968
rect 5718 8956 5724 8968
rect 5679 8928 5724 8956
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 6472 8965 6500 9132
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 7653 9027 7711 9033
rect 7653 9024 7665 9027
rect 6696 8996 7665 9024
rect 6696 8984 6702 8996
rect 7653 8993 7665 8996
rect 7699 8993 7711 9027
rect 7653 8987 7711 8993
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 1854 8848 1860 8900
rect 1912 8888 1918 8900
rect 2961 8891 3019 8897
rect 2961 8888 2973 8891
rect 1912 8860 2973 8888
rect 1912 8848 1918 8860
rect 2961 8857 2973 8860
rect 3007 8857 3019 8891
rect 2961 8851 3019 8857
rect 5476 8891 5534 8897
rect 5476 8857 5488 8891
rect 5522 8888 5534 8891
rect 5522 8860 7144 8888
rect 5522 8857 5534 8860
rect 5476 8851 5534 8857
rect 1946 8820 1952 8832
rect 1907 8792 1952 8820
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 2866 8820 2872 8832
rect 2827 8792 2872 8820
rect 2866 8780 2872 8792
rect 2924 8780 2930 8832
rect 4154 8780 4160 8832
rect 4212 8820 4218 8832
rect 4341 8823 4399 8829
rect 4341 8820 4353 8823
rect 4212 8792 4353 8820
rect 4212 8780 4218 8792
rect 4341 8789 4353 8792
rect 4387 8789 4399 8823
rect 4341 8783 4399 8789
rect 6641 8823 6699 8829
rect 6641 8789 6653 8823
rect 6687 8820 6699 8823
rect 6822 8820 6828 8832
rect 6687 8792 6828 8820
rect 6687 8789 6699 8792
rect 6641 8783 6699 8789
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 7116 8829 7144 8860
rect 7101 8823 7159 8829
rect 7101 8789 7113 8823
rect 7147 8789 7159 8823
rect 7466 8820 7472 8832
rect 7427 8792 7472 8820
rect 7101 8783 7159 8789
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 7558 8780 7564 8832
rect 7616 8820 7622 8832
rect 7616 8792 7661 8820
rect 7616 8780 7622 8792
rect 1104 8730 8556 8752
rect 1104 8678 3466 8730
rect 3518 8678 3530 8730
rect 3582 8678 3594 8730
rect 3646 8678 3658 8730
rect 3710 8678 5950 8730
rect 6002 8678 6014 8730
rect 6066 8678 6078 8730
rect 6130 8678 6142 8730
rect 6194 8678 8556 8730
rect 1104 8656 8556 8678
rect 2317 8619 2375 8625
rect 2317 8585 2329 8619
rect 2363 8616 2375 8619
rect 2866 8616 2872 8628
rect 2363 8588 2872 8616
rect 2363 8585 2375 8588
rect 2317 8579 2375 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 5718 8616 5724 8628
rect 4448 8588 5724 8616
rect 14 8508 20 8560
rect 72 8548 78 8560
rect 1581 8551 1639 8557
rect 1581 8548 1593 8551
rect 72 8520 1593 8548
rect 72 8508 78 8520
rect 1581 8517 1593 8520
rect 1627 8517 1639 8551
rect 1581 8511 1639 8517
rect 1765 8551 1823 8557
rect 1765 8517 1777 8551
rect 1811 8548 1823 8551
rect 1854 8548 1860 8560
rect 1811 8520 1860 8548
rect 1811 8517 1823 8520
rect 1765 8511 1823 8517
rect 1854 8508 1860 8520
rect 1912 8508 1918 8560
rect 3441 8483 3499 8489
rect 3441 8449 3453 8483
rect 3487 8480 3499 8483
rect 3786 8480 3792 8492
rect 3487 8452 3792 8480
rect 3487 8449 3499 8452
rect 3441 8443 3499 8449
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 4448 8489 4476 8588
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 6365 8619 6423 8625
rect 6365 8585 6377 8619
rect 6411 8585 6423 8619
rect 6822 8616 6828 8628
rect 6783 8588 6828 8616
rect 6365 8579 6423 8585
rect 4700 8551 4758 8557
rect 4700 8517 4712 8551
rect 4746 8548 4758 8551
rect 6380 8548 6408 8579
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 4746 8520 6408 8548
rect 4746 8517 4758 8520
rect 4700 8511 4758 8517
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8449 4491 8483
rect 4433 8443 4491 8449
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 6733 8483 6791 8489
rect 6733 8480 6745 8483
rect 5592 8452 6745 8480
rect 5592 8440 5598 8452
rect 6733 8449 6745 8452
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8480 7895 8483
rect 8294 8480 8300 8492
rect 7883 8452 8300 8480
rect 7883 8449 7895 8452
rect 7837 8443 7895 8449
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 3694 8412 3700 8424
rect 3655 8384 3700 8412
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 6638 8372 6644 8424
rect 6696 8412 6702 8424
rect 6822 8412 6828 8424
rect 6696 8384 6828 8412
rect 6696 8372 6702 8384
rect 6822 8372 6828 8384
rect 6880 8412 6886 8424
rect 6917 8415 6975 8421
rect 6917 8412 6929 8415
rect 6880 8384 6929 8412
rect 6880 8372 6886 8384
rect 6917 8381 6929 8384
rect 6963 8381 6975 8415
rect 6917 8375 6975 8381
rect 5813 8347 5871 8353
rect 5813 8313 5825 8347
rect 5859 8344 5871 8347
rect 7466 8344 7472 8356
rect 5859 8316 7472 8344
rect 5859 8313 5871 8316
rect 5813 8307 5871 8313
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 7650 8276 7656 8288
rect 7611 8248 7656 8276
rect 7650 8236 7656 8248
rect 7708 8236 7714 8288
rect 1104 8186 8556 8208
rect 1104 8134 2224 8186
rect 2276 8134 2288 8186
rect 2340 8134 2352 8186
rect 2404 8134 2416 8186
rect 2468 8134 4708 8186
rect 4760 8134 4772 8186
rect 4824 8134 4836 8186
rect 4888 8134 4900 8186
rect 4952 8134 7192 8186
rect 7244 8134 7256 8186
rect 7308 8134 7320 8186
rect 7372 8134 7384 8186
rect 7436 8134 8556 8186
rect 1104 8112 8556 8134
rect 1854 8072 1860 8084
rect 1815 8044 1860 8072
rect 1854 8032 1860 8044
rect 1912 8032 1918 8084
rect 3786 8072 3792 8084
rect 3747 8044 3792 8072
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 6549 8075 6607 8081
rect 6549 8072 6561 8075
rect 5776 8044 6561 8072
rect 5776 8032 5782 8044
rect 6549 8041 6561 8044
rect 6595 8041 6607 8075
rect 6549 8035 6607 8041
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 7616 8044 7665 8072
rect 7616 8032 7622 8044
rect 7653 8041 7665 8044
rect 7699 8041 7711 8075
rect 7653 8035 7711 8041
rect 3237 7939 3295 7945
rect 3237 7905 3249 7939
rect 3283 7936 3295 7939
rect 3326 7936 3332 7948
rect 3283 7908 3332 7936
rect 3283 7905 3295 7908
rect 3237 7899 3295 7905
rect 3326 7896 3332 7908
rect 3384 7936 3390 7948
rect 3694 7936 3700 7948
rect 3384 7908 3700 7936
rect 3384 7896 3390 7908
rect 3694 7896 3700 7908
rect 3752 7896 3758 7948
rect 4338 7936 4344 7948
rect 4299 7908 4344 7936
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 2958 7828 2964 7880
rect 3016 7877 3022 7880
rect 3016 7868 3028 7877
rect 4154 7868 4160 7880
rect 3016 7840 3061 7868
rect 4115 7840 4160 7868
rect 3016 7831 3028 7840
rect 3016 7828 3022 7831
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 6788 7840 7849 7868
rect 6788 7828 6794 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 5258 7800 5264 7812
rect 5219 7772 5264 7800
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 4246 7692 4252 7744
rect 4304 7732 4310 7744
rect 4304 7704 4349 7732
rect 4304 7692 4310 7704
rect 1104 7642 8556 7664
rect 1104 7590 3466 7642
rect 3518 7590 3530 7642
rect 3582 7590 3594 7642
rect 3646 7590 3658 7642
rect 3710 7590 5950 7642
rect 6002 7590 6014 7642
rect 6066 7590 6078 7642
rect 6130 7590 6142 7642
rect 6194 7590 8556 7642
rect 1104 7568 8556 7590
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 5353 7531 5411 7537
rect 5353 7528 5365 7531
rect 5316 7500 5365 7528
rect 5316 7488 5322 7500
rect 5353 7497 5365 7500
rect 5399 7497 5411 7531
rect 5353 7491 5411 7497
rect 6365 7531 6423 7537
rect 6365 7497 6377 7531
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 6825 7531 6883 7537
rect 6825 7497 6837 7531
rect 6871 7528 6883 7531
rect 7650 7528 7656 7540
rect 6871 7500 7656 7528
rect 6871 7497 6883 7500
rect 6825 7491 6883 7497
rect 2308 7463 2366 7469
rect 2308 7429 2320 7463
rect 2354 7460 2366 7463
rect 6380 7460 6408 7491
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 2354 7432 6408 7460
rect 2354 7429 2366 7432
rect 2308 7423 2366 7429
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7392 2099 7395
rect 3326 7392 3332 7404
rect 2087 7364 3332 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 4065 7395 4123 7401
rect 4065 7361 4077 7395
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 7006 7392 7012 7404
rect 6779 7364 7012 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 3050 7284 3056 7336
rect 3108 7324 3114 7336
rect 4080 7324 4108 7355
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 3108 7296 4108 7324
rect 6840 7296 6929 7324
rect 3108 7284 3114 7296
rect 6840 7200 6868 7296
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 3421 7191 3479 7197
rect 3421 7188 3433 7191
rect 3292 7160 3433 7188
rect 3292 7148 3298 7160
rect 3421 7157 3433 7160
rect 3467 7157 3479 7191
rect 3421 7151 3479 7157
rect 4338 7148 4344 7200
rect 4396 7188 4402 7200
rect 6822 7188 6828 7200
rect 4396 7160 6828 7188
rect 4396 7148 4402 7160
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 1104 7098 8556 7120
rect 1104 7046 2224 7098
rect 2276 7046 2288 7098
rect 2340 7046 2352 7098
rect 2404 7046 2416 7098
rect 2468 7046 4708 7098
rect 4760 7046 4772 7098
rect 4824 7046 4836 7098
rect 4888 7046 4900 7098
rect 4952 7046 7192 7098
rect 7244 7046 7256 7098
rect 7308 7046 7320 7098
rect 7372 7046 7384 7098
rect 7436 7046 8556 7098
rect 1104 7024 8556 7046
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7101 6987 7159 6993
rect 7101 6984 7113 6987
rect 7064 6956 7113 6984
rect 7064 6944 7070 6956
rect 7101 6953 7113 6956
rect 7147 6953 7159 6987
rect 7101 6947 7159 6953
rect 5718 6848 5724 6860
rect 5679 6820 5724 6848
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 3237 6783 3295 6789
rect 3237 6780 3249 6783
rect 3200 6752 3249 6780
rect 3200 6740 3206 6752
rect 3237 6749 3249 6752
rect 3283 6780 3295 6783
rect 3326 6780 3332 6792
rect 3283 6752 3332 6780
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 3881 6783 3939 6789
rect 3881 6749 3893 6783
rect 3927 6780 3939 6783
rect 5736 6780 5764 6808
rect 3927 6752 5764 6780
rect 3927 6749 3939 6752
rect 3881 6743 3939 6749
rect 2866 6672 2872 6724
rect 2924 6712 2930 6724
rect 2970 6715 3028 6721
rect 2970 6712 2982 6715
rect 2924 6684 2982 6712
rect 2924 6672 2930 6684
rect 2970 6681 2982 6684
rect 3016 6681 3028 6715
rect 2970 6675 3028 6681
rect 4148 6715 4206 6721
rect 4148 6681 4160 6715
rect 4194 6712 4206 6715
rect 5442 6712 5448 6724
rect 4194 6684 5448 6712
rect 4194 6681 4206 6684
rect 4148 6675 4206 6681
rect 5442 6672 5448 6684
rect 5500 6672 5506 6724
rect 5988 6715 6046 6721
rect 5988 6681 6000 6715
rect 6034 6712 6046 6715
rect 6362 6712 6368 6724
rect 6034 6684 6368 6712
rect 6034 6681 6046 6684
rect 5988 6675 6046 6681
rect 6362 6672 6368 6684
rect 6420 6672 6426 6724
rect 1854 6644 1860 6656
rect 1815 6616 1860 6644
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5534 6644 5540 6656
rect 5307 6616 5540 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 1104 6554 8556 6576
rect 1104 6502 3466 6554
rect 3518 6502 3530 6554
rect 3582 6502 3594 6554
rect 3646 6502 3658 6554
rect 3710 6502 5950 6554
rect 6002 6502 6014 6554
rect 6066 6502 6078 6554
rect 6130 6502 6142 6554
rect 6194 6502 8556 6554
rect 1104 6480 8556 6502
rect 2866 6440 2872 6452
rect 2827 6412 2872 6440
rect 2866 6400 2872 6412
rect 2924 6400 2930 6452
rect 3234 6440 3240 6452
rect 3195 6412 3240 6440
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 5442 6400 5448 6452
rect 5500 6440 5506 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 5500 6412 6377 6440
rect 5500 6400 5506 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 1946 6332 1952 6384
rect 2004 6372 2010 6384
rect 3329 6375 3387 6381
rect 3329 6372 3341 6375
rect 2004 6344 3341 6372
rect 2004 6332 2010 6344
rect 3329 6341 3341 6344
rect 3375 6341 3387 6375
rect 5718 6372 5724 6384
rect 3329 6335 3387 6341
rect 4448 6344 5724 6372
rect 4448 6313 4476 6344
rect 5718 6332 5724 6344
rect 5776 6332 5782 6384
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6273 4491 6307
rect 4433 6267 4491 6273
rect 4700 6307 4758 6313
rect 4700 6273 4712 6307
rect 4746 6304 4758 6307
rect 5074 6304 5080 6316
rect 4746 6276 5080 6304
rect 4746 6273 4758 6276
rect 4700 6267 4758 6273
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 5166 6264 5172 6316
rect 5224 6304 5230 6316
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 5224 6276 6745 6304
rect 5224 6264 5230 6276
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 7834 6304 7840 6316
rect 7795 6276 7840 6304
rect 6733 6267 6791 6273
rect 7834 6264 7840 6276
rect 7892 6264 7898 6316
rect 3513 6239 3571 6245
rect 3513 6205 3525 6239
rect 3559 6236 3571 6239
rect 4338 6236 4344 6248
rect 3559 6208 4344 6236
rect 3559 6205 3571 6208
rect 3513 6199 3571 6205
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 6822 6236 6828 6248
rect 6783 6208 6828 6236
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 7006 6236 7012 6248
rect 6967 6208 7012 6236
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 5813 6103 5871 6109
rect 5813 6069 5825 6103
rect 5859 6100 5871 6103
rect 5994 6100 6000 6112
rect 5859 6072 6000 6100
rect 5859 6069 5871 6072
rect 5813 6063 5871 6069
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 6270 6060 6276 6112
rect 6328 6100 6334 6112
rect 7653 6103 7711 6109
rect 7653 6100 7665 6103
rect 6328 6072 7665 6100
rect 6328 6060 6334 6072
rect 7653 6069 7665 6072
rect 7699 6069 7711 6103
rect 7653 6063 7711 6069
rect 1104 6010 8556 6032
rect 1104 5958 2224 6010
rect 2276 5958 2288 6010
rect 2340 5958 2352 6010
rect 2404 5958 2416 6010
rect 2468 5958 4708 6010
rect 4760 5958 4772 6010
rect 4824 5958 4836 6010
rect 4888 5958 4900 6010
rect 4952 5958 7192 6010
rect 7244 5958 7256 6010
rect 7308 5958 7320 6010
rect 7372 5958 7384 6010
rect 7436 5958 8556 6010
rect 1104 5936 8556 5958
rect 5166 5896 5172 5908
rect 5127 5868 5172 5896
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 6362 5896 6368 5908
rect 6323 5868 6368 5896
rect 6362 5856 6368 5868
rect 6420 5856 6426 5908
rect 5813 5763 5871 5769
rect 5813 5729 5825 5763
rect 5859 5760 5871 5763
rect 7006 5760 7012 5772
rect 5859 5732 7012 5760
rect 5859 5729 5871 5732
rect 5813 5723 5871 5729
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 3142 5692 3148 5704
rect 2884 5664 3148 5692
rect 2884 5568 2912 5664
rect 3142 5652 3148 5664
rect 3200 5692 3206 5704
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3200 5664 3801 5692
rect 3200 5652 3206 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 5350 5692 5356 5704
rect 3789 5655 3847 5661
rect 3988 5664 5356 5692
rect 3237 5627 3295 5633
rect 3237 5593 3249 5627
rect 3283 5624 3295 5627
rect 3988 5624 4016 5664
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 5994 5692 6000 5704
rect 5955 5664 6000 5692
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 3283 5596 4016 5624
rect 4056 5627 4114 5633
rect 3283 5593 3295 5596
rect 3237 5587 3295 5593
rect 4056 5593 4068 5627
rect 4102 5624 4114 5627
rect 4706 5624 4712 5636
rect 4102 5596 4712 5624
rect 4102 5593 4114 5596
rect 4056 5587 4114 5593
rect 4706 5584 4712 5596
rect 4764 5584 4770 5636
rect 1949 5559 2007 5565
rect 1949 5525 1961 5559
rect 1995 5556 2007 5559
rect 2866 5556 2872 5568
rect 1995 5528 2872 5556
rect 1995 5525 2007 5528
rect 1949 5519 2007 5525
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 5905 5559 5963 5565
rect 5905 5556 5917 5559
rect 5684 5528 5917 5556
rect 5684 5516 5690 5528
rect 5905 5525 5917 5528
rect 5951 5525 5963 5559
rect 5905 5519 5963 5525
rect 1104 5466 8556 5488
rect 1104 5414 3466 5466
rect 3518 5414 3530 5466
rect 3582 5414 3594 5466
rect 3646 5414 3658 5466
rect 3710 5414 5950 5466
rect 6002 5414 6014 5466
rect 6066 5414 6078 5466
rect 6130 5414 6142 5466
rect 6194 5414 8556 5466
rect 1104 5392 8556 5414
rect 1854 5312 1860 5364
rect 1912 5352 1918 5364
rect 2041 5355 2099 5361
rect 2041 5352 2053 5355
rect 1912 5324 2053 5352
rect 1912 5312 1918 5324
rect 2041 5321 2053 5324
rect 2087 5321 2099 5355
rect 2041 5315 2099 5321
rect 2409 5355 2467 5361
rect 2409 5321 2421 5355
rect 2455 5321 2467 5355
rect 2409 5315 2467 5321
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 5077 5355 5135 5361
rect 5077 5352 5089 5355
rect 4295 5324 5089 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 5077 5321 5089 5324
rect 5123 5321 5135 5355
rect 5077 5315 5135 5321
rect 2424 5284 2452 5315
rect 3114 5287 3172 5293
rect 3114 5284 3126 5287
rect 2424 5256 3126 5284
rect 3114 5253 3126 5256
rect 3160 5253 3172 5287
rect 3114 5247 3172 5253
rect 5169 5219 5227 5225
rect 1780 5188 4844 5216
rect 1780 5157 1808 5188
rect 1765 5151 1823 5157
rect 1765 5117 1777 5151
rect 1811 5117 1823 5151
rect 1946 5148 1952 5160
rect 1907 5120 1952 5148
rect 1765 5111 1823 5117
rect 1946 5108 1952 5120
rect 2004 5108 2010 5160
rect 2866 5148 2872 5160
rect 2827 5120 2872 5148
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 4816 5148 4844 5188
rect 5169 5185 5181 5219
rect 5215 5216 5227 5219
rect 7650 5216 7656 5228
rect 5215 5188 7656 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 5258 5148 5264 5160
rect 4816 5120 5264 5148
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 4706 5080 4712 5092
rect 4667 5052 4712 5080
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 1104 4922 8556 4944
rect 1104 4870 2224 4922
rect 2276 4870 2288 4922
rect 2340 4870 2352 4922
rect 2404 4870 2416 4922
rect 2468 4870 4708 4922
rect 4760 4870 4772 4922
rect 4824 4870 4836 4922
rect 4888 4870 4900 4922
rect 4952 4870 7192 4922
rect 7244 4870 7256 4922
rect 7308 4870 7320 4922
rect 7372 4870 7384 4922
rect 7436 4870 8556 4922
rect 1104 4848 8556 4870
rect 4985 4811 5043 4817
rect 4985 4777 4997 4811
rect 5031 4808 5043 4811
rect 5074 4808 5080 4820
rect 5031 4780 5080 4808
rect 5031 4777 5043 4780
rect 4985 4771 5043 4777
rect 5074 4768 5080 4780
rect 5132 4768 5138 4820
rect 6270 4672 6276 4684
rect 5184 4644 6276 4672
rect 5184 4613 5212 4644
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 7006 4604 7012 4616
rect 5316 4576 7012 4604
rect 5316 4564 5322 4576
rect 7006 4564 7012 4576
rect 7064 4564 7070 4616
rect 1104 4378 8556 4400
rect 1104 4326 3466 4378
rect 3518 4326 3530 4378
rect 3582 4326 3594 4378
rect 3646 4326 3658 4378
rect 3710 4326 5950 4378
rect 6002 4326 6014 4378
rect 6066 4326 6078 4378
rect 6130 4326 6142 4378
rect 6194 4326 8556 4378
rect 1104 4304 8556 4326
rect 1762 4128 1768 4140
rect 1723 4100 1768 4128
rect 1762 4088 1768 4100
rect 1820 4088 1826 4140
rect 1949 3995 2007 4001
rect 1949 3961 1961 3995
rect 1995 3992 2007 3995
rect 6822 3992 6828 4004
rect 1995 3964 6828 3992
rect 1995 3961 2007 3964
rect 1949 3955 2007 3961
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 1104 3834 8556 3856
rect 1104 3782 2224 3834
rect 2276 3782 2288 3834
rect 2340 3782 2352 3834
rect 2404 3782 2416 3834
rect 2468 3782 4708 3834
rect 4760 3782 4772 3834
rect 4824 3782 4836 3834
rect 4888 3782 4900 3834
rect 4952 3782 7192 3834
rect 7244 3782 7256 3834
rect 7308 3782 7320 3834
rect 7372 3782 7384 3834
rect 7436 3782 8556 3834
rect 1104 3760 8556 3782
rect 1104 3290 8556 3312
rect 1104 3238 3466 3290
rect 3518 3238 3530 3290
rect 3582 3238 3594 3290
rect 3646 3238 3658 3290
rect 3710 3238 5950 3290
rect 6002 3238 6014 3290
rect 6066 3238 6078 3290
rect 6130 3238 6142 3290
rect 6194 3238 8556 3290
rect 1104 3216 8556 3238
rect 7650 3176 7656 3188
rect 7611 3148 7656 3176
rect 7650 3136 7656 3148
rect 7708 3136 7714 3188
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 8110 3040 8116 3052
rect 7883 3012 8116 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 1104 2746 8556 2768
rect 1104 2694 2224 2746
rect 2276 2694 2288 2746
rect 2340 2694 2352 2746
rect 2404 2694 2416 2746
rect 2468 2694 4708 2746
rect 4760 2694 4772 2746
rect 4824 2694 4836 2746
rect 4888 2694 4900 2746
rect 4952 2694 7192 2746
rect 7244 2694 7256 2746
rect 7308 2694 7320 2746
rect 7372 2694 7384 2746
rect 7436 2694 8556 2746
rect 1104 2672 8556 2694
rect 1946 2632 1952 2644
rect 1907 2604 1952 2632
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 4246 2632 4252 2644
rect 2915 2604 4252 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 5626 2632 5632 2644
rect 5587 2604 5632 2632
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 7469 2635 7527 2641
rect 7469 2632 7481 2635
rect 7064 2604 7481 2632
rect 7064 2592 7070 2604
rect 7469 2601 7481 2604
rect 7515 2601 7527 2635
rect 7469 2595 7527 2601
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 72 2400 1777 2428
rect 72 2388 78 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2590 2388 2596 2440
rect 2648 2428 2654 2440
rect 2685 2431 2743 2437
rect 2685 2428 2697 2431
rect 2648 2400 2697 2428
rect 2648 2388 2654 2400
rect 2685 2397 2697 2400
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 5350 2388 5356 2440
rect 5408 2428 5414 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5408 2400 5457 2428
rect 5408 2388 5414 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 7742 2360 7748 2372
rect 7703 2332 7748 2360
rect 7742 2320 7748 2332
rect 7800 2320 7806 2372
rect 1104 2202 8556 2224
rect 1104 2150 3466 2202
rect 3518 2150 3530 2202
rect 3582 2150 3594 2202
rect 3646 2150 3658 2202
rect 3710 2150 5950 2202
rect 6002 2150 6014 2202
rect 6066 2150 6078 2202
rect 6130 2150 6142 2202
rect 6194 2150 8556 2202
rect 1104 2128 8556 2150
<< via1 >>
rect 2224 9222 2276 9274
rect 2288 9222 2340 9274
rect 2352 9222 2404 9274
rect 2416 9222 2468 9274
rect 4708 9222 4760 9274
rect 4772 9222 4824 9274
rect 4836 9222 4888 9274
rect 4900 9222 4952 9274
rect 7192 9222 7244 9274
rect 7256 9222 7308 9274
rect 7320 9222 7372 9274
rect 7384 9222 7436 9274
rect 5540 9120 5592 9172
rect 2964 9052 3016 9104
rect 4344 8984 4396 9036
rect 1768 8959 1820 8968
rect 1768 8925 1777 8959
rect 1777 8925 1811 8959
rect 1811 8925 1820 8959
rect 1768 8916 1820 8925
rect 5724 8959 5776 8968
rect 5724 8925 5733 8959
rect 5733 8925 5767 8959
rect 5767 8925 5776 8959
rect 5724 8916 5776 8925
rect 6644 8984 6696 9036
rect 1860 8848 1912 8900
rect 1952 8823 2004 8832
rect 1952 8789 1961 8823
rect 1961 8789 1995 8823
rect 1995 8789 2004 8823
rect 1952 8780 2004 8789
rect 2872 8823 2924 8832
rect 2872 8789 2881 8823
rect 2881 8789 2915 8823
rect 2915 8789 2924 8823
rect 2872 8780 2924 8789
rect 4160 8780 4212 8832
rect 6828 8780 6880 8832
rect 7472 8823 7524 8832
rect 7472 8789 7481 8823
rect 7481 8789 7515 8823
rect 7515 8789 7524 8823
rect 7472 8780 7524 8789
rect 7564 8823 7616 8832
rect 7564 8789 7573 8823
rect 7573 8789 7607 8823
rect 7607 8789 7616 8823
rect 7564 8780 7616 8789
rect 3466 8678 3518 8730
rect 3530 8678 3582 8730
rect 3594 8678 3646 8730
rect 3658 8678 3710 8730
rect 5950 8678 6002 8730
rect 6014 8678 6066 8730
rect 6078 8678 6130 8730
rect 6142 8678 6194 8730
rect 2872 8576 2924 8628
rect 20 8508 72 8560
rect 1860 8508 1912 8560
rect 3792 8440 3844 8492
rect 5724 8576 5776 8628
rect 6828 8619 6880 8628
rect 6828 8585 6837 8619
rect 6837 8585 6871 8619
rect 6871 8585 6880 8619
rect 6828 8576 6880 8585
rect 5540 8440 5592 8492
rect 8300 8440 8352 8492
rect 3700 8415 3752 8424
rect 3700 8381 3709 8415
rect 3709 8381 3743 8415
rect 3743 8381 3752 8415
rect 3700 8372 3752 8381
rect 6644 8372 6696 8424
rect 6828 8372 6880 8424
rect 7472 8304 7524 8356
rect 7656 8279 7708 8288
rect 7656 8245 7665 8279
rect 7665 8245 7699 8279
rect 7699 8245 7708 8279
rect 7656 8236 7708 8245
rect 2224 8134 2276 8186
rect 2288 8134 2340 8186
rect 2352 8134 2404 8186
rect 2416 8134 2468 8186
rect 4708 8134 4760 8186
rect 4772 8134 4824 8186
rect 4836 8134 4888 8186
rect 4900 8134 4952 8186
rect 7192 8134 7244 8186
rect 7256 8134 7308 8186
rect 7320 8134 7372 8186
rect 7384 8134 7436 8186
rect 1860 8075 1912 8084
rect 1860 8041 1869 8075
rect 1869 8041 1903 8075
rect 1903 8041 1912 8075
rect 1860 8032 1912 8041
rect 3792 8075 3844 8084
rect 3792 8041 3801 8075
rect 3801 8041 3835 8075
rect 3835 8041 3844 8075
rect 3792 8032 3844 8041
rect 5724 8032 5776 8084
rect 7564 8032 7616 8084
rect 3332 7896 3384 7948
rect 3700 7896 3752 7948
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 2964 7871 3016 7880
rect 2964 7837 2982 7871
rect 2982 7837 3016 7871
rect 4160 7871 4212 7880
rect 2964 7828 3016 7837
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 6736 7828 6788 7880
rect 5264 7803 5316 7812
rect 5264 7769 5273 7803
rect 5273 7769 5307 7803
rect 5307 7769 5316 7803
rect 5264 7760 5316 7769
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 3466 7590 3518 7642
rect 3530 7590 3582 7642
rect 3594 7590 3646 7642
rect 3658 7590 3710 7642
rect 5950 7590 6002 7642
rect 6014 7590 6066 7642
rect 6078 7590 6130 7642
rect 6142 7590 6194 7642
rect 5264 7488 5316 7540
rect 7656 7488 7708 7540
rect 3332 7352 3384 7404
rect 3056 7284 3108 7336
rect 7012 7352 7064 7404
rect 3240 7148 3292 7200
rect 4344 7148 4396 7200
rect 6828 7148 6880 7200
rect 2224 7046 2276 7098
rect 2288 7046 2340 7098
rect 2352 7046 2404 7098
rect 2416 7046 2468 7098
rect 4708 7046 4760 7098
rect 4772 7046 4824 7098
rect 4836 7046 4888 7098
rect 4900 7046 4952 7098
rect 7192 7046 7244 7098
rect 7256 7046 7308 7098
rect 7320 7046 7372 7098
rect 7384 7046 7436 7098
rect 7012 6944 7064 6996
rect 5724 6851 5776 6860
rect 5724 6817 5733 6851
rect 5733 6817 5767 6851
rect 5767 6817 5776 6851
rect 5724 6808 5776 6817
rect 3148 6740 3200 6792
rect 3332 6740 3384 6792
rect 2872 6672 2924 6724
rect 5448 6672 5500 6724
rect 6368 6672 6420 6724
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 5540 6604 5592 6656
rect 3466 6502 3518 6554
rect 3530 6502 3582 6554
rect 3594 6502 3646 6554
rect 3658 6502 3710 6554
rect 5950 6502 6002 6554
rect 6014 6502 6066 6554
rect 6078 6502 6130 6554
rect 6142 6502 6194 6554
rect 2872 6443 2924 6452
rect 2872 6409 2881 6443
rect 2881 6409 2915 6443
rect 2915 6409 2924 6443
rect 2872 6400 2924 6409
rect 3240 6443 3292 6452
rect 3240 6409 3249 6443
rect 3249 6409 3283 6443
rect 3283 6409 3292 6443
rect 3240 6400 3292 6409
rect 5448 6400 5500 6452
rect 1952 6332 2004 6384
rect 5724 6332 5776 6384
rect 5080 6264 5132 6316
rect 5172 6264 5224 6316
rect 7840 6307 7892 6316
rect 7840 6273 7849 6307
rect 7849 6273 7883 6307
rect 7883 6273 7892 6307
rect 7840 6264 7892 6273
rect 4344 6196 4396 6248
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 7012 6239 7064 6248
rect 7012 6205 7021 6239
rect 7021 6205 7055 6239
rect 7055 6205 7064 6239
rect 7012 6196 7064 6205
rect 6000 6060 6052 6112
rect 6276 6060 6328 6112
rect 2224 5958 2276 6010
rect 2288 5958 2340 6010
rect 2352 5958 2404 6010
rect 2416 5958 2468 6010
rect 4708 5958 4760 6010
rect 4772 5958 4824 6010
rect 4836 5958 4888 6010
rect 4900 5958 4952 6010
rect 7192 5958 7244 6010
rect 7256 5958 7308 6010
rect 7320 5958 7372 6010
rect 7384 5958 7436 6010
rect 5172 5899 5224 5908
rect 5172 5865 5181 5899
rect 5181 5865 5215 5899
rect 5215 5865 5224 5899
rect 5172 5856 5224 5865
rect 6368 5899 6420 5908
rect 6368 5865 6377 5899
rect 6377 5865 6411 5899
rect 6411 5865 6420 5899
rect 6368 5856 6420 5865
rect 7012 5720 7064 5772
rect 3148 5652 3200 5704
rect 5356 5652 5408 5704
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 4712 5584 4764 5636
rect 2872 5516 2924 5568
rect 5632 5516 5684 5568
rect 3466 5414 3518 5466
rect 3530 5414 3582 5466
rect 3594 5414 3646 5466
rect 3658 5414 3710 5466
rect 5950 5414 6002 5466
rect 6014 5414 6066 5466
rect 6078 5414 6130 5466
rect 6142 5414 6194 5466
rect 1860 5312 1912 5364
rect 1952 5151 2004 5160
rect 1952 5117 1961 5151
rect 1961 5117 1995 5151
rect 1995 5117 2004 5151
rect 1952 5108 2004 5117
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 7656 5176 7708 5228
rect 5264 5151 5316 5160
rect 5264 5117 5273 5151
rect 5273 5117 5307 5151
rect 5307 5117 5316 5151
rect 5264 5108 5316 5117
rect 4712 5083 4764 5092
rect 4712 5049 4721 5083
rect 4721 5049 4755 5083
rect 4755 5049 4764 5083
rect 4712 5040 4764 5049
rect 2224 4870 2276 4922
rect 2288 4870 2340 4922
rect 2352 4870 2404 4922
rect 2416 4870 2468 4922
rect 4708 4870 4760 4922
rect 4772 4870 4824 4922
rect 4836 4870 4888 4922
rect 4900 4870 4952 4922
rect 7192 4870 7244 4922
rect 7256 4870 7308 4922
rect 7320 4870 7372 4922
rect 7384 4870 7436 4922
rect 5080 4768 5132 4820
rect 6276 4632 6328 4684
rect 5264 4607 5316 4616
rect 5264 4573 5273 4607
rect 5273 4573 5307 4607
rect 5307 4573 5316 4607
rect 5264 4564 5316 4573
rect 7012 4564 7064 4616
rect 3466 4326 3518 4378
rect 3530 4326 3582 4378
rect 3594 4326 3646 4378
rect 3658 4326 3710 4378
rect 5950 4326 6002 4378
rect 6014 4326 6066 4378
rect 6078 4326 6130 4378
rect 6142 4326 6194 4378
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 6828 3952 6880 4004
rect 2224 3782 2276 3834
rect 2288 3782 2340 3834
rect 2352 3782 2404 3834
rect 2416 3782 2468 3834
rect 4708 3782 4760 3834
rect 4772 3782 4824 3834
rect 4836 3782 4888 3834
rect 4900 3782 4952 3834
rect 7192 3782 7244 3834
rect 7256 3782 7308 3834
rect 7320 3782 7372 3834
rect 7384 3782 7436 3834
rect 3466 3238 3518 3290
rect 3530 3238 3582 3290
rect 3594 3238 3646 3290
rect 3658 3238 3710 3290
rect 5950 3238 6002 3290
rect 6014 3238 6066 3290
rect 6078 3238 6130 3290
rect 6142 3238 6194 3290
rect 7656 3179 7708 3188
rect 7656 3145 7665 3179
rect 7665 3145 7699 3179
rect 7699 3145 7708 3179
rect 7656 3136 7708 3145
rect 8116 3000 8168 3052
rect 2224 2694 2276 2746
rect 2288 2694 2340 2746
rect 2352 2694 2404 2746
rect 2416 2694 2468 2746
rect 4708 2694 4760 2746
rect 4772 2694 4824 2746
rect 4836 2694 4888 2746
rect 4900 2694 4952 2746
rect 7192 2694 7244 2746
rect 7256 2694 7308 2746
rect 7320 2694 7372 2746
rect 7384 2694 7436 2746
rect 1952 2635 2004 2644
rect 1952 2601 1961 2635
rect 1961 2601 1995 2635
rect 1995 2601 2004 2635
rect 1952 2592 2004 2601
rect 4252 2592 4304 2644
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 7012 2592 7064 2644
rect 20 2388 72 2440
rect 2596 2388 2648 2440
rect 5356 2388 5408 2440
rect 7748 2363 7800 2372
rect 7748 2329 7757 2363
rect 7757 2329 7791 2363
rect 7791 2329 7800 2363
rect 7748 2320 7800 2329
rect 3466 2150 3518 2202
rect 3530 2150 3582 2202
rect 3594 2150 3646 2202
rect 3658 2150 3710 2202
rect 5950 2150 6002 2202
rect 6014 2150 6066 2202
rect 6078 2150 6130 2202
rect 6142 2150 6194 2202
<< metal2 >>
rect 18 11079 74 11879
rect 2778 11079 2834 11879
rect 32 8566 60 11079
rect 2792 10962 2820 11079
rect 2884 11070 3096 11098
rect 5538 11079 5594 11879
rect 8298 11079 8354 11879
rect 2884 10962 2912 11070
rect 2792 10934 2912 10962
rect 2198 9276 2494 9296
rect 2254 9274 2278 9276
rect 2334 9274 2358 9276
rect 2414 9274 2438 9276
rect 2276 9222 2278 9274
rect 2340 9222 2352 9274
rect 2414 9222 2416 9274
rect 2254 9220 2278 9222
rect 2334 9220 2358 9222
rect 2414 9220 2438 9222
rect 2198 9200 2494 9220
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 20 8560 72 8566
rect 20 8502 72 8508
rect 1780 7993 1808 8910
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 8566 1900 8842
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 1860 8560 1912 8566
rect 1860 8502 1912 8508
rect 1872 8090 1900 8502
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1766 7984 1822 7993
rect 1766 7919 1822 7928
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 5370 1900 6598
rect 1964 6390 1992 8774
rect 2884 8634 2912 8774
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2198 8188 2494 8208
rect 2254 8186 2278 8188
rect 2334 8186 2358 8188
rect 2414 8186 2438 8188
rect 2276 8134 2278 8186
rect 2340 8134 2352 8186
rect 2414 8134 2416 8186
rect 2254 8132 2278 8134
rect 2334 8132 2358 8134
rect 2414 8132 2438 8134
rect 2198 8112 2494 8132
rect 2976 7886 3004 9046
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 3068 7342 3096 11070
rect 4682 9276 4978 9296
rect 4738 9274 4762 9276
rect 4818 9274 4842 9276
rect 4898 9274 4922 9276
rect 4760 9222 4762 9274
rect 4824 9222 4836 9274
rect 4898 9222 4900 9274
rect 4738 9220 4762 9222
rect 4818 9220 4842 9222
rect 4898 9220 4922 9222
rect 4682 9200 4978 9220
rect 5552 9178 5580 11079
rect 6734 9888 6790 9897
rect 6734 9823 6790 9832
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 3440 8732 3736 8752
rect 3496 8730 3520 8732
rect 3576 8730 3600 8732
rect 3656 8730 3680 8732
rect 3518 8678 3520 8730
rect 3582 8678 3594 8730
rect 3656 8678 3658 8730
rect 3496 8676 3520 8678
rect 3576 8676 3600 8678
rect 3656 8676 3680 8678
rect 3440 8656 3736 8676
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3712 7954 3740 8366
rect 3804 8090 3832 8434
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3344 7410 3372 7890
rect 4172 7886 4200 8774
rect 4356 7954 4384 8978
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5736 8634 5764 8910
rect 5924 8732 6220 8752
rect 5980 8730 6004 8732
rect 6060 8730 6084 8732
rect 6140 8730 6164 8732
rect 6002 8678 6004 8730
rect 6066 8678 6078 8730
rect 6140 8678 6142 8730
rect 5980 8676 6004 8678
rect 6060 8676 6084 8678
rect 6140 8676 6164 8678
rect 5924 8656 6220 8676
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 4682 8188 4978 8208
rect 4738 8186 4762 8188
rect 4818 8186 4842 8188
rect 4898 8186 4922 8188
rect 4760 8134 4762 8186
rect 4824 8134 4836 8186
rect 4898 8134 4900 8186
rect 4738 8132 4762 8134
rect 4818 8132 4842 8134
rect 4898 8132 4922 8134
rect 4682 8112 4978 8132
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 3440 7644 3736 7664
rect 3496 7642 3520 7644
rect 3576 7642 3600 7644
rect 3656 7642 3680 7644
rect 3518 7590 3520 7642
rect 3582 7590 3594 7642
rect 3656 7590 3658 7642
rect 3496 7588 3520 7590
rect 3576 7588 3600 7590
rect 3656 7588 3680 7590
rect 3440 7568 3736 7588
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 2198 7100 2494 7120
rect 2254 7098 2278 7100
rect 2334 7098 2358 7100
rect 2414 7098 2438 7100
rect 2276 7046 2278 7098
rect 2340 7046 2352 7098
rect 2414 7046 2416 7098
rect 2254 7044 2278 7046
rect 2334 7044 2358 7046
rect 2414 7044 2438 7046
rect 2198 7024 2494 7044
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2884 6458 2912 6666
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 1952 6384 2004 6390
rect 1952 6326 2004 6332
rect 2198 6012 2494 6032
rect 2254 6010 2278 6012
rect 2334 6010 2358 6012
rect 2414 6010 2438 6012
rect 2276 5958 2278 6010
rect 2340 5958 2352 6010
rect 2414 5958 2416 6010
rect 2254 5956 2278 5958
rect 2334 5956 2358 5958
rect 2414 5956 2438 5958
rect 2198 5936 2494 5956
rect 3160 5710 3188 6734
rect 3252 6458 3280 7142
rect 3344 6798 3372 7346
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3440 6556 3736 6576
rect 3496 6554 3520 6556
rect 3576 6554 3600 6556
rect 3656 6554 3680 6556
rect 3518 6502 3520 6554
rect 3582 6502 3594 6554
rect 3656 6502 3658 6554
rect 3496 6500 3520 6502
rect 3576 6500 3600 6502
rect 3656 6500 3680 6502
rect 3440 6480 3736 6500
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 2884 5166 2912 5510
rect 3440 5468 3736 5488
rect 3496 5466 3520 5468
rect 3576 5466 3600 5468
rect 3656 5466 3680 5468
rect 3518 5414 3520 5466
rect 3582 5414 3594 5466
rect 3656 5414 3658 5466
rect 3496 5412 3520 5414
rect 3576 5412 3600 5414
rect 3656 5412 3680 5414
rect 3440 5392 3736 5412
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1780 3913 1808 4082
rect 1766 3904 1822 3913
rect 1766 3839 1822 3848
rect 1964 2650 1992 5102
rect 2198 4924 2494 4944
rect 2254 4922 2278 4924
rect 2334 4922 2358 4924
rect 2414 4922 2438 4924
rect 2276 4870 2278 4922
rect 2340 4870 2352 4922
rect 2414 4870 2416 4922
rect 2254 4868 2278 4870
rect 2334 4868 2358 4870
rect 2414 4868 2438 4870
rect 2198 4848 2494 4868
rect 3440 4380 3736 4400
rect 3496 4378 3520 4380
rect 3576 4378 3600 4380
rect 3656 4378 3680 4380
rect 3518 4326 3520 4378
rect 3582 4326 3594 4378
rect 3656 4326 3658 4378
rect 3496 4324 3520 4326
rect 3576 4324 3600 4326
rect 3656 4324 3680 4326
rect 3440 4304 3736 4324
rect 2198 3836 2494 3856
rect 2254 3834 2278 3836
rect 2334 3834 2358 3836
rect 2414 3834 2438 3836
rect 2276 3782 2278 3834
rect 2340 3782 2352 3834
rect 2414 3782 2416 3834
rect 2254 3780 2278 3782
rect 2334 3780 2358 3782
rect 2414 3780 2438 3782
rect 2198 3760 2494 3780
rect 3440 3292 3736 3312
rect 3496 3290 3520 3292
rect 3576 3290 3600 3292
rect 3656 3290 3680 3292
rect 3518 3238 3520 3290
rect 3582 3238 3594 3290
rect 3656 3238 3658 3290
rect 3496 3236 3520 3238
rect 3576 3236 3600 3238
rect 3656 3236 3680 3238
rect 3440 3216 3736 3236
rect 2198 2748 2494 2768
rect 2254 2746 2278 2748
rect 2334 2746 2358 2748
rect 2414 2746 2438 2748
rect 2276 2694 2278 2746
rect 2340 2694 2352 2746
rect 2414 2694 2416 2746
rect 2254 2692 2278 2694
rect 2334 2692 2358 2694
rect 2414 2692 2438 2694
rect 2198 2672 2494 2692
rect 4264 2650 4292 7686
rect 4356 7206 4384 7890
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5276 7546 5304 7754
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4356 6254 4384 7142
rect 4682 7100 4978 7120
rect 4738 7098 4762 7100
rect 4818 7098 4842 7100
rect 4898 7098 4922 7100
rect 4760 7046 4762 7098
rect 4824 7046 4836 7098
rect 4898 7046 4900 7098
rect 4738 7044 4762 7046
rect 4818 7044 4842 7046
rect 4898 7044 4922 7046
rect 4682 7024 4978 7044
rect 5276 6914 5304 7482
rect 5276 6886 5396 6914
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4682 6012 4978 6032
rect 4738 6010 4762 6012
rect 4818 6010 4842 6012
rect 4898 6010 4922 6012
rect 4760 5958 4762 6010
rect 4824 5958 4836 6010
rect 4898 5958 4900 6010
rect 4738 5956 4762 5958
rect 4818 5956 4842 5958
rect 4898 5956 4922 5958
rect 4682 5936 4978 5956
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4724 5098 4752 5578
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4682 4924 4978 4944
rect 4738 4922 4762 4924
rect 4818 4922 4842 4924
rect 4898 4922 4922 4924
rect 4760 4870 4762 4922
rect 4824 4870 4836 4922
rect 4898 4870 4900 4922
rect 4738 4868 4762 4870
rect 4818 4868 4842 4870
rect 4898 4868 4922 4870
rect 4682 4848 4978 4868
rect 5092 4826 5120 6258
rect 5184 5914 5212 6258
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5368 5710 5396 6886
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5460 6458 5488 6666
rect 5552 6662 5580 8434
rect 5736 8090 5764 8570
rect 6656 8430 6684 8978
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5736 6866 5764 8026
rect 6748 7886 6776 9823
rect 7166 9276 7462 9296
rect 7222 9274 7246 9276
rect 7302 9274 7326 9276
rect 7382 9274 7406 9276
rect 7244 9222 7246 9274
rect 7308 9222 7320 9274
rect 7382 9222 7384 9274
rect 7222 9220 7246 9222
rect 7302 9220 7326 9222
rect 7382 9220 7406 9222
rect 7166 9200 7462 9220
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 6840 8634 6868 8774
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 5924 7644 6220 7664
rect 5980 7642 6004 7644
rect 6060 7642 6084 7644
rect 6140 7642 6164 7644
rect 6002 7590 6004 7642
rect 6066 7590 6078 7642
rect 6140 7590 6142 7642
rect 5980 7588 6004 7590
rect 6060 7588 6084 7590
rect 6140 7588 6164 7590
rect 5924 7568 6220 7588
rect 6840 7206 6868 8366
rect 7484 8362 7512 8774
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7166 8188 7462 8208
rect 7222 8186 7246 8188
rect 7302 8186 7326 8188
rect 7382 8186 7406 8188
rect 7244 8134 7246 8186
rect 7308 8134 7320 8186
rect 7382 8134 7384 8186
rect 7222 8132 7246 8134
rect 7302 8132 7326 8134
rect 7382 8132 7406 8134
rect 7166 8112 7462 8132
rect 7576 8090 7604 8774
rect 8312 8498 8340 11079
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7668 7546 7696 8230
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5736 6390 5764 6802
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 5924 6556 6220 6576
rect 5980 6554 6004 6556
rect 6060 6554 6084 6556
rect 6140 6554 6164 6556
rect 6002 6502 6004 6554
rect 6066 6502 6078 6554
rect 6140 6502 6142 6554
rect 5980 6500 6004 6502
rect 6060 6500 6084 6502
rect 6140 6500 6164 6502
rect 5924 6480 6220 6500
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6012 5710 6040 6054
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5276 4622 5304 5102
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 4682 3836 4978 3856
rect 4738 3834 4762 3836
rect 4818 3834 4842 3836
rect 4898 3834 4922 3836
rect 4760 3782 4762 3834
rect 4824 3782 4836 3834
rect 4898 3782 4900 3834
rect 4738 3780 4762 3782
rect 4818 3780 4842 3782
rect 4898 3780 4922 3782
rect 4682 3760 4978 3780
rect 4682 2748 4978 2768
rect 4738 2746 4762 2748
rect 4818 2746 4842 2748
rect 4898 2746 4922 2748
rect 4760 2694 4762 2746
rect 4824 2694 4836 2746
rect 4898 2694 4900 2746
rect 4738 2692 4762 2694
rect 4818 2692 4842 2694
rect 4898 2692 4922 2694
rect 4682 2672 4978 2692
rect 5644 2650 5672 5510
rect 5924 5468 6220 5488
rect 5980 5466 6004 5468
rect 6060 5466 6084 5468
rect 6140 5466 6164 5468
rect 6002 5414 6004 5466
rect 6066 5414 6078 5466
rect 6140 5414 6142 5466
rect 5980 5412 6004 5414
rect 6060 5412 6084 5414
rect 6140 5412 6164 5414
rect 5924 5392 6220 5412
rect 6288 4690 6316 6054
rect 6380 5914 6408 6666
rect 6840 6338 6868 7142
rect 7024 7002 7052 7346
rect 7166 7100 7462 7120
rect 7222 7098 7246 7100
rect 7302 7098 7326 7100
rect 7382 7098 7406 7100
rect 7244 7046 7246 7098
rect 7308 7046 7320 7098
rect 7382 7046 7384 7098
rect 7222 7044 7246 7046
rect 7302 7044 7326 7046
rect 7382 7044 7406 7046
rect 7166 7024 7462 7044
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6840 6310 7052 6338
rect 7024 6254 7052 6310
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 5924 4380 6220 4400
rect 5980 4378 6004 4380
rect 6060 4378 6084 4380
rect 6140 4378 6164 4380
rect 6002 4326 6004 4378
rect 6066 4326 6078 4378
rect 6140 4326 6142 4378
rect 5980 4324 6004 4326
rect 6060 4324 6084 4326
rect 6140 4324 6164 4326
rect 5924 4304 6220 4324
rect 6840 4010 6868 6190
rect 7024 5778 7052 6190
rect 7166 6012 7462 6032
rect 7222 6010 7246 6012
rect 7302 6010 7326 6012
rect 7382 6010 7406 6012
rect 7244 5958 7246 6010
rect 7308 5958 7320 6010
rect 7382 5958 7384 6010
rect 7222 5956 7246 5958
rect 7302 5956 7326 5958
rect 7382 5956 7406 5958
rect 7166 5936 7462 5956
rect 7852 5817 7880 6258
rect 7838 5808 7894 5817
rect 7012 5772 7064 5778
rect 7838 5743 7894 5752
rect 7012 5714 7064 5720
rect 7024 4622 7052 5714
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7166 4924 7462 4944
rect 7222 4922 7246 4924
rect 7302 4922 7326 4924
rect 7382 4922 7406 4924
rect 7244 4870 7246 4922
rect 7308 4870 7320 4922
rect 7382 4870 7384 4922
rect 7222 4868 7246 4870
rect 7302 4868 7326 4870
rect 7382 4868 7406 4870
rect 7166 4848 7462 4868
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 5924 3292 6220 3312
rect 5980 3290 6004 3292
rect 6060 3290 6084 3292
rect 6140 3290 6164 3292
rect 6002 3238 6004 3290
rect 6066 3238 6078 3290
rect 6140 3238 6142 3290
rect 5980 3236 6004 3238
rect 6060 3236 6084 3238
rect 6140 3236 6164 3238
rect 5924 3216 6220 3236
rect 7024 2650 7052 4558
rect 7166 3836 7462 3856
rect 7222 3834 7246 3836
rect 7302 3834 7326 3836
rect 7382 3834 7406 3836
rect 7244 3782 7246 3834
rect 7308 3782 7320 3834
rect 7382 3782 7384 3834
rect 7222 3780 7246 3782
rect 7302 3780 7326 3782
rect 7382 3780 7406 3782
rect 7166 3760 7462 3780
rect 7668 3194 7696 5170
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 7166 2748 7462 2768
rect 7222 2746 7246 2748
rect 7302 2746 7326 2748
rect 7382 2746 7406 2748
rect 7244 2694 7246 2746
rect 7308 2694 7320 2746
rect 7382 2694 7384 2746
rect 7222 2692 7246 2694
rect 7302 2692 7326 2694
rect 7382 2692 7406 2694
rect 7166 2672 7462 2692
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 32 800 60 2382
rect 2608 800 2636 2382
rect 3440 2204 3736 2224
rect 3496 2202 3520 2204
rect 3576 2202 3600 2204
rect 3656 2202 3680 2204
rect 3518 2150 3520 2202
rect 3582 2150 3594 2202
rect 3656 2150 3658 2202
rect 3496 2148 3520 2150
rect 3576 2148 3600 2150
rect 3656 2148 3680 2150
rect 3440 2128 3736 2148
rect 5368 800 5396 2382
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 5924 2204 6220 2224
rect 5980 2202 6004 2204
rect 6060 2202 6084 2204
rect 6140 2202 6164 2204
rect 6002 2150 6004 2202
rect 6066 2150 6078 2202
rect 6140 2150 6142 2202
rect 5980 2148 6004 2150
rect 6060 2148 6084 2150
rect 6140 2148 6164 2150
rect 5924 2128 6220 2148
rect 7760 1737 7788 2314
rect 7746 1728 7802 1737
rect 7746 1663 7802 1672
rect 8128 800 8156 2994
rect 18 0 74 800
rect 2594 0 2650 800
rect 5354 0 5410 800
rect 8114 0 8170 800
<< via2 >>
rect 2198 9274 2254 9276
rect 2278 9274 2334 9276
rect 2358 9274 2414 9276
rect 2438 9274 2494 9276
rect 2198 9222 2224 9274
rect 2224 9222 2254 9274
rect 2278 9222 2288 9274
rect 2288 9222 2334 9274
rect 2358 9222 2404 9274
rect 2404 9222 2414 9274
rect 2438 9222 2468 9274
rect 2468 9222 2494 9274
rect 2198 9220 2254 9222
rect 2278 9220 2334 9222
rect 2358 9220 2414 9222
rect 2438 9220 2494 9222
rect 1766 7928 1822 7984
rect 2198 8186 2254 8188
rect 2278 8186 2334 8188
rect 2358 8186 2414 8188
rect 2438 8186 2494 8188
rect 2198 8134 2224 8186
rect 2224 8134 2254 8186
rect 2278 8134 2288 8186
rect 2288 8134 2334 8186
rect 2358 8134 2404 8186
rect 2404 8134 2414 8186
rect 2438 8134 2468 8186
rect 2468 8134 2494 8186
rect 2198 8132 2254 8134
rect 2278 8132 2334 8134
rect 2358 8132 2414 8134
rect 2438 8132 2494 8134
rect 4682 9274 4738 9276
rect 4762 9274 4818 9276
rect 4842 9274 4898 9276
rect 4922 9274 4978 9276
rect 4682 9222 4708 9274
rect 4708 9222 4738 9274
rect 4762 9222 4772 9274
rect 4772 9222 4818 9274
rect 4842 9222 4888 9274
rect 4888 9222 4898 9274
rect 4922 9222 4952 9274
rect 4952 9222 4978 9274
rect 4682 9220 4738 9222
rect 4762 9220 4818 9222
rect 4842 9220 4898 9222
rect 4922 9220 4978 9222
rect 6734 9832 6790 9888
rect 3440 8730 3496 8732
rect 3520 8730 3576 8732
rect 3600 8730 3656 8732
rect 3680 8730 3736 8732
rect 3440 8678 3466 8730
rect 3466 8678 3496 8730
rect 3520 8678 3530 8730
rect 3530 8678 3576 8730
rect 3600 8678 3646 8730
rect 3646 8678 3656 8730
rect 3680 8678 3710 8730
rect 3710 8678 3736 8730
rect 3440 8676 3496 8678
rect 3520 8676 3576 8678
rect 3600 8676 3656 8678
rect 3680 8676 3736 8678
rect 5924 8730 5980 8732
rect 6004 8730 6060 8732
rect 6084 8730 6140 8732
rect 6164 8730 6220 8732
rect 5924 8678 5950 8730
rect 5950 8678 5980 8730
rect 6004 8678 6014 8730
rect 6014 8678 6060 8730
rect 6084 8678 6130 8730
rect 6130 8678 6140 8730
rect 6164 8678 6194 8730
rect 6194 8678 6220 8730
rect 5924 8676 5980 8678
rect 6004 8676 6060 8678
rect 6084 8676 6140 8678
rect 6164 8676 6220 8678
rect 4682 8186 4738 8188
rect 4762 8186 4818 8188
rect 4842 8186 4898 8188
rect 4922 8186 4978 8188
rect 4682 8134 4708 8186
rect 4708 8134 4738 8186
rect 4762 8134 4772 8186
rect 4772 8134 4818 8186
rect 4842 8134 4888 8186
rect 4888 8134 4898 8186
rect 4922 8134 4952 8186
rect 4952 8134 4978 8186
rect 4682 8132 4738 8134
rect 4762 8132 4818 8134
rect 4842 8132 4898 8134
rect 4922 8132 4978 8134
rect 3440 7642 3496 7644
rect 3520 7642 3576 7644
rect 3600 7642 3656 7644
rect 3680 7642 3736 7644
rect 3440 7590 3466 7642
rect 3466 7590 3496 7642
rect 3520 7590 3530 7642
rect 3530 7590 3576 7642
rect 3600 7590 3646 7642
rect 3646 7590 3656 7642
rect 3680 7590 3710 7642
rect 3710 7590 3736 7642
rect 3440 7588 3496 7590
rect 3520 7588 3576 7590
rect 3600 7588 3656 7590
rect 3680 7588 3736 7590
rect 2198 7098 2254 7100
rect 2278 7098 2334 7100
rect 2358 7098 2414 7100
rect 2438 7098 2494 7100
rect 2198 7046 2224 7098
rect 2224 7046 2254 7098
rect 2278 7046 2288 7098
rect 2288 7046 2334 7098
rect 2358 7046 2404 7098
rect 2404 7046 2414 7098
rect 2438 7046 2468 7098
rect 2468 7046 2494 7098
rect 2198 7044 2254 7046
rect 2278 7044 2334 7046
rect 2358 7044 2414 7046
rect 2438 7044 2494 7046
rect 2198 6010 2254 6012
rect 2278 6010 2334 6012
rect 2358 6010 2414 6012
rect 2438 6010 2494 6012
rect 2198 5958 2224 6010
rect 2224 5958 2254 6010
rect 2278 5958 2288 6010
rect 2288 5958 2334 6010
rect 2358 5958 2404 6010
rect 2404 5958 2414 6010
rect 2438 5958 2468 6010
rect 2468 5958 2494 6010
rect 2198 5956 2254 5958
rect 2278 5956 2334 5958
rect 2358 5956 2414 5958
rect 2438 5956 2494 5958
rect 3440 6554 3496 6556
rect 3520 6554 3576 6556
rect 3600 6554 3656 6556
rect 3680 6554 3736 6556
rect 3440 6502 3466 6554
rect 3466 6502 3496 6554
rect 3520 6502 3530 6554
rect 3530 6502 3576 6554
rect 3600 6502 3646 6554
rect 3646 6502 3656 6554
rect 3680 6502 3710 6554
rect 3710 6502 3736 6554
rect 3440 6500 3496 6502
rect 3520 6500 3576 6502
rect 3600 6500 3656 6502
rect 3680 6500 3736 6502
rect 3440 5466 3496 5468
rect 3520 5466 3576 5468
rect 3600 5466 3656 5468
rect 3680 5466 3736 5468
rect 3440 5414 3466 5466
rect 3466 5414 3496 5466
rect 3520 5414 3530 5466
rect 3530 5414 3576 5466
rect 3600 5414 3646 5466
rect 3646 5414 3656 5466
rect 3680 5414 3710 5466
rect 3710 5414 3736 5466
rect 3440 5412 3496 5414
rect 3520 5412 3576 5414
rect 3600 5412 3656 5414
rect 3680 5412 3736 5414
rect 1766 3848 1822 3904
rect 2198 4922 2254 4924
rect 2278 4922 2334 4924
rect 2358 4922 2414 4924
rect 2438 4922 2494 4924
rect 2198 4870 2224 4922
rect 2224 4870 2254 4922
rect 2278 4870 2288 4922
rect 2288 4870 2334 4922
rect 2358 4870 2404 4922
rect 2404 4870 2414 4922
rect 2438 4870 2468 4922
rect 2468 4870 2494 4922
rect 2198 4868 2254 4870
rect 2278 4868 2334 4870
rect 2358 4868 2414 4870
rect 2438 4868 2494 4870
rect 3440 4378 3496 4380
rect 3520 4378 3576 4380
rect 3600 4378 3656 4380
rect 3680 4378 3736 4380
rect 3440 4326 3466 4378
rect 3466 4326 3496 4378
rect 3520 4326 3530 4378
rect 3530 4326 3576 4378
rect 3600 4326 3646 4378
rect 3646 4326 3656 4378
rect 3680 4326 3710 4378
rect 3710 4326 3736 4378
rect 3440 4324 3496 4326
rect 3520 4324 3576 4326
rect 3600 4324 3656 4326
rect 3680 4324 3736 4326
rect 2198 3834 2254 3836
rect 2278 3834 2334 3836
rect 2358 3834 2414 3836
rect 2438 3834 2494 3836
rect 2198 3782 2224 3834
rect 2224 3782 2254 3834
rect 2278 3782 2288 3834
rect 2288 3782 2334 3834
rect 2358 3782 2404 3834
rect 2404 3782 2414 3834
rect 2438 3782 2468 3834
rect 2468 3782 2494 3834
rect 2198 3780 2254 3782
rect 2278 3780 2334 3782
rect 2358 3780 2414 3782
rect 2438 3780 2494 3782
rect 3440 3290 3496 3292
rect 3520 3290 3576 3292
rect 3600 3290 3656 3292
rect 3680 3290 3736 3292
rect 3440 3238 3466 3290
rect 3466 3238 3496 3290
rect 3520 3238 3530 3290
rect 3530 3238 3576 3290
rect 3600 3238 3646 3290
rect 3646 3238 3656 3290
rect 3680 3238 3710 3290
rect 3710 3238 3736 3290
rect 3440 3236 3496 3238
rect 3520 3236 3576 3238
rect 3600 3236 3656 3238
rect 3680 3236 3736 3238
rect 2198 2746 2254 2748
rect 2278 2746 2334 2748
rect 2358 2746 2414 2748
rect 2438 2746 2494 2748
rect 2198 2694 2224 2746
rect 2224 2694 2254 2746
rect 2278 2694 2288 2746
rect 2288 2694 2334 2746
rect 2358 2694 2404 2746
rect 2404 2694 2414 2746
rect 2438 2694 2468 2746
rect 2468 2694 2494 2746
rect 2198 2692 2254 2694
rect 2278 2692 2334 2694
rect 2358 2692 2414 2694
rect 2438 2692 2494 2694
rect 4682 7098 4738 7100
rect 4762 7098 4818 7100
rect 4842 7098 4898 7100
rect 4922 7098 4978 7100
rect 4682 7046 4708 7098
rect 4708 7046 4738 7098
rect 4762 7046 4772 7098
rect 4772 7046 4818 7098
rect 4842 7046 4888 7098
rect 4888 7046 4898 7098
rect 4922 7046 4952 7098
rect 4952 7046 4978 7098
rect 4682 7044 4738 7046
rect 4762 7044 4818 7046
rect 4842 7044 4898 7046
rect 4922 7044 4978 7046
rect 4682 6010 4738 6012
rect 4762 6010 4818 6012
rect 4842 6010 4898 6012
rect 4922 6010 4978 6012
rect 4682 5958 4708 6010
rect 4708 5958 4738 6010
rect 4762 5958 4772 6010
rect 4772 5958 4818 6010
rect 4842 5958 4888 6010
rect 4888 5958 4898 6010
rect 4922 5958 4952 6010
rect 4952 5958 4978 6010
rect 4682 5956 4738 5958
rect 4762 5956 4818 5958
rect 4842 5956 4898 5958
rect 4922 5956 4978 5958
rect 4682 4922 4738 4924
rect 4762 4922 4818 4924
rect 4842 4922 4898 4924
rect 4922 4922 4978 4924
rect 4682 4870 4708 4922
rect 4708 4870 4738 4922
rect 4762 4870 4772 4922
rect 4772 4870 4818 4922
rect 4842 4870 4888 4922
rect 4888 4870 4898 4922
rect 4922 4870 4952 4922
rect 4952 4870 4978 4922
rect 4682 4868 4738 4870
rect 4762 4868 4818 4870
rect 4842 4868 4898 4870
rect 4922 4868 4978 4870
rect 7166 9274 7222 9276
rect 7246 9274 7302 9276
rect 7326 9274 7382 9276
rect 7406 9274 7462 9276
rect 7166 9222 7192 9274
rect 7192 9222 7222 9274
rect 7246 9222 7256 9274
rect 7256 9222 7302 9274
rect 7326 9222 7372 9274
rect 7372 9222 7382 9274
rect 7406 9222 7436 9274
rect 7436 9222 7462 9274
rect 7166 9220 7222 9222
rect 7246 9220 7302 9222
rect 7326 9220 7382 9222
rect 7406 9220 7462 9222
rect 5924 7642 5980 7644
rect 6004 7642 6060 7644
rect 6084 7642 6140 7644
rect 6164 7642 6220 7644
rect 5924 7590 5950 7642
rect 5950 7590 5980 7642
rect 6004 7590 6014 7642
rect 6014 7590 6060 7642
rect 6084 7590 6130 7642
rect 6130 7590 6140 7642
rect 6164 7590 6194 7642
rect 6194 7590 6220 7642
rect 5924 7588 5980 7590
rect 6004 7588 6060 7590
rect 6084 7588 6140 7590
rect 6164 7588 6220 7590
rect 7166 8186 7222 8188
rect 7246 8186 7302 8188
rect 7326 8186 7382 8188
rect 7406 8186 7462 8188
rect 7166 8134 7192 8186
rect 7192 8134 7222 8186
rect 7246 8134 7256 8186
rect 7256 8134 7302 8186
rect 7326 8134 7372 8186
rect 7372 8134 7382 8186
rect 7406 8134 7436 8186
rect 7436 8134 7462 8186
rect 7166 8132 7222 8134
rect 7246 8132 7302 8134
rect 7326 8132 7382 8134
rect 7406 8132 7462 8134
rect 5924 6554 5980 6556
rect 6004 6554 6060 6556
rect 6084 6554 6140 6556
rect 6164 6554 6220 6556
rect 5924 6502 5950 6554
rect 5950 6502 5980 6554
rect 6004 6502 6014 6554
rect 6014 6502 6060 6554
rect 6084 6502 6130 6554
rect 6130 6502 6140 6554
rect 6164 6502 6194 6554
rect 6194 6502 6220 6554
rect 5924 6500 5980 6502
rect 6004 6500 6060 6502
rect 6084 6500 6140 6502
rect 6164 6500 6220 6502
rect 4682 3834 4738 3836
rect 4762 3834 4818 3836
rect 4842 3834 4898 3836
rect 4922 3834 4978 3836
rect 4682 3782 4708 3834
rect 4708 3782 4738 3834
rect 4762 3782 4772 3834
rect 4772 3782 4818 3834
rect 4842 3782 4888 3834
rect 4888 3782 4898 3834
rect 4922 3782 4952 3834
rect 4952 3782 4978 3834
rect 4682 3780 4738 3782
rect 4762 3780 4818 3782
rect 4842 3780 4898 3782
rect 4922 3780 4978 3782
rect 4682 2746 4738 2748
rect 4762 2746 4818 2748
rect 4842 2746 4898 2748
rect 4922 2746 4978 2748
rect 4682 2694 4708 2746
rect 4708 2694 4738 2746
rect 4762 2694 4772 2746
rect 4772 2694 4818 2746
rect 4842 2694 4888 2746
rect 4888 2694 4898 2746
rect 4922 2694 4952 2746
rect 4952 2694 4978 2746
rect 4682 2692 4738 2694
rect 4762 2692 4818 2694
rect 4842 2692 4898 2694
rect 4922 2692 4978 2694
rect 5924 5466 5980 5468
rect 6004 5466 6060 5468
rect 6084 5466 6140 5468
rect 6164 5466 6220 5468
rect 5924 5414 5950 5466
rect 5950 5414 5980 5466
rect 6004 5414 6014 5466
rect 6014 5414 6060 5466
rect 6084 5414 6130 5466
rect 6130 5414 6140 5466
rect 6164 5414 6194 5466
rect 6194 5414 6220 5466
rect 5924 5412 5980 5414
rect 6004 5412 6060 5414
rect 6084 5412 6140 5414
rect 6164 5412 6220 5414
rect 7166 7098 7222 7100
rect 7246 7098 7302 7100
rect 7326 7098 7382 7100
rect 7406 7098 7462 7100
rect 7166 7046 7192 7098
rect 7192 7046 7222 7098
rect 7246 7046 7256 7098
rect 7256 7046 7302 7098
rect 7326 7046 7372 7098
rect 7372 7046 7382 7098
rect 7406 7046 7436 7098
rect 7436 7046 7462 7098
rect 7166 7044 7222 7046
rect 7246 7044 7302 7046
rect 7326 7044 7382 7046
rect 7406 7044 7462 7046
rect 5924 4378 5980 4380
rect 6004 4378 6060 4380
rect 6084 4378 6140 4380
rect 6164 4378 6220 4380
rect 5924 4326 5950 4378
rect 5950 4326 5980 4378
rect 6004 4326 6014 4378
rect 6014 4326 6060 4378
rect 6084 4326 6130 4378
rect 6130 4326 6140 4378
rect 6164 4326 6194 4378
rect 6194 4326 6220 4378
rect 5924 4324 5980 4326
rect 6004 4324 6060 4326
rect 6084 4324 6140 4326
rect 6164 4324 6220 4326
rect 7166 6010 7222 6012
rect 7246 6010 7302 6012
rect 7326 6010 7382 6012
rect 7406 6010 7462 6012
rect 7166 5958 7192 6010
rect 7192 5958 7222 6010
rect 7246 5958 7256 6010
rect 7256 5958 7302 6010
rect 7326 5958 7372 6010
rect 7372 5958 7382 6010
rect 7406 5958 7436 6010
rect 7436 5958 7462 6010
rect 7166 5956 7222 5958
rect 7246 5956 7302 5958
rect 7326 5956 7382 5958
rect 7406 5956 7462 5958
rect 7838 5752 7894 5808
rect 7166 4922 7222 4924
rect 7246 4922 7302 4924
rect 7326 4922 7382 4924
rect 7406 4922 7462 4924
rect 7166 4870 7192 4922
rect 7192 4870 7222 4922
rect 7246 4870 7256 4922
rect 7256 4870 7302 4922
rect 7326 4870 7372 4922
rect 7372 4870 7382 4922
rect 7406 4870 7436 4922
rect 7436 4870 7462 4922
rect 7166 4868 7222 4870
rect 7246 4868 7302 4870
rect 7326 4868 7382 4870
rect 7406 4868 7462 4870
rect 5924 3290 5980 3292
rect 6004 3290 6060 3292
rect 6084 3290 6140 3292
rect 6164 3290 6220 3292
rect 5924 3238 5950 3290
rect 5950 3238 5980 3290
rect 6004 3238 6014 3290
rect 6014 3238 6060 3290
rect 6084 3238 6130 3290
rect 6130 3238 6140 3290
rect 6164 3238 6194 3290
rect 6194 3238 6220 3290
rect 5924 3236 5980 3238
rect 6004 3236 6060 3238
rect 6084 3236 6140 3238
rect 6164 3236 6220 3238
rect 7166 3834 7222 3836
rect 7246 3834 7302 3836
rect 7326 3834 7382 3836
rect 7406 3834 7462 3836
rect 7166 3782 7192 3834
rect 7192 3782 7222 3834
rect 7246 3782 7256 3834
rect 7256 3782 7302 3834
rect 7326 3782 7372 3834
rect 7372 3782 7382 3834
rect 7406 3782 7436 3834
rect 7436 3782 7462 3834
rect 7166 3780 7222 3782
rect 7246 3780 7302 3782
rect 7326 3780 7382 3782
rect 7406 3780 7462 3782
rect 7166 2746 7222 2748
rect 7246 2746 7302 2748
rect 7326 2746 7382 2748
rect 7406 2746 7462 2748
rect 7166 2694 7192 2746
rect 7192 2694 7222 2746
rect 7246 2694 7256 2746
rect 7256 2694 7302 2746
rect 7326 2694 7372 2746
rect 7372 2694 7382 2746
rect 7406 2694 7436 2746
rect 7436 2694 7462 2746
rect 7166 2692 7222 2694
rect 7246 2692 7302 2694
rect 7326 2692 7382 2694
rect 7406 2692 7462 2694
rect 3440 2202 3496 2204
rect 3520 2202 3576 2204
rect 3600 2202 3656 2204
rect 3680 2202 3736 2204
rect 3440 2150 3466 2202
rect 3466 2150 3496 2202
rect 3520 2150 3530 2202
rect 3530 2150 3576 2202
rect 3600 2150 3646 2202
rect 3646 2150 3656 2202
rect 3680 2150 3710 2202
rect 3710 2150 3736 2202
rect 3440 2148 3496 2150
rect 3520 2148 3576 2150
rect 3600 2148 3656 2150
rect 3680 2148 3736 2150
rect 5924 2202 5980 2204
rect 6004 2202 6060 2204
rect 6084 2202 6140 2204
rect 6164 2202 6220 2204
rect 5924 2150 5950 2202
rect 5950 2150 5980 2202
rect 6004 2150 6014 2202
rect 6014 2150 6060 2202
rect 6084 2150 6130 2202
rect 6130 2150 6140 2202
rect 6164 2150 6194 2202
rect 6194 2150 6220 2202
rect 5924 2148 5980 2150
rect 6004 2148 6060 2150
rect 6084 2148 6140 2150
rect 6164 2148 6220 2150
rect 7746 1672 7802 1728
<< metal3 >>
rect 6729 9890 6795 9893
rect 8935 9890 9735 9920
rect 6729 9888 9735 9890
rect 6729 9832 6734 9888
rect 6790 9832 9735 9888
rect 6729 9830 9735 9832
rect 6729 9827 6795 9830
rect 8935 9800 9735 9830
rect 2186 9280 2506 9281
rect 2186 9216 2194 9280
rect 2258 9216 2274 9280
rect 2338 9216 2354 9280
rect 2418 9216 2434 9280
rect 2498 9216 2506 9280
rect 2186 9215 2506 9216
rect 4670 9280 4990 9281
rect 4670 9216 4678 9280
rect 4742 9216 4758 9280
rect 4822 9216 4838 9280
rect 4902 9216 4918 9280
rect 4982 9216 4990 9280
rect 4670 9215 4990 9216
rect 7154 9280 7474 9281
rect 7154 9216 7162 9280
rect 7226 9216 7242 9280
rect 7306 9216 7322 9280
rect 7386 9216 7402 9280
rect 7466 9216 7474 9280
rect 7154 9215 7474 9216
rect 3428 8736 3748 8737
rect 3428 8672 3436 8736
rect 3500 8672 3516 8736
rect 3580 8672 3596 8736
rect 3660 8672 3676 8736
rect 3740 8672 3748 8736
rect 3428 8671 3748 8672
rect 5912 8736 6232 8737
rect 5912 8672 5920 8736
rect 5984 8672 6000 8736
rect 6064 8672 6080 8736
rect 6144 8672 6160 8736
rect 6224 8672 6232 8736
rect 5912 8671 6232 8672
rect 2186 8192 2506 8193
rect 2186 8128 2194 8192
rect 2258 8128 2274 8192
rect 2338 8128 2354 8192
rect 2418 8128 2434 8192
rect 2498 8128 2506 8192
rect 2186 8127 2506 8128
rect 4670 8192 4990 8193
rect 4670 8128 4678 8192
rect 4742 8128 4758 8192
rect 4822 8128 4838 8192
rect 4902 8128 4918 8192
rect 4982 8128 4990 8192
rect 4670 8127 4990 8128
rect 7154 8192 7474 8193
rect 7154 8128 7162 8192
rect 7226 8128 7242 8192
rect 7306 8128 7322 8192
rect 7386 8128 7402 8192
rect 7466 8128 7474 8192
rect 7154 8127 7474 8128
rect 0 7986 800 8016
rect 1761 7986 1827 7989
rect 0 7984 1827 7986
rect 0 7928 1766 7984
rect 1822 7928 1827 7984
rect 0 7926 1827 7928
rect 0 7896 800 7926
rect 1761 7923 1827 7926
rect 3428 7648 3748 7649
rect 3428 7584 3436 7648
rect 3500 7584 3516 7648
rect 3580 7584 3596 7648
rect 3660 7584 3676 7648
rect 3740 7584 3748 7648
rect 3428 7583 3748 7584
rect 5912 7648 6232 7649
rect 5912 7584 5920 7648
rect 5984 7584 6000 7648
rect 6064 7584 6080 7648
rect 6144 7584 6160 7648
rect 6224 7584 6232 7648
rect 5912 7583 6232 7584
rect 2186 7104 2506 7105
rect 2186 7040 2194 7104
rect 2258 7040 2274 7104
rect 2338 7040 2354 7104
rect 2418 7040 2434 7104
rect 2498 7040 2506 7104
rect 2186 7039 2506 7040
rect 4670 7104 4990 7105
rect 4670 7040 4678 7104
rect 4742 7040 4758 7104
rect 4822 7040 4838 7104
rect 4902 7040 4918 7104
rect 4982 7040 4990 7104
rect 4670 7039 4990 7040
rect 7154 7104 7474 7105
rect 7154 7040 7162 7104
rect 7226 7040 7242 7104
rect 7306 7040 7322 7104
rect 7386 7040 7402 7104
rect 7466 7040 7474 7104
rect 7154 7039 7474 7040
rect 3428 6560 3748 6561
rect 3428 6496 3436 6560
rect 3500 6496 3516 6560
rect 3580 6496 3596 6560
rect 3660 6496 3676 6560
rect 3740 6496 3748 6560
rect 3428 6495 3748 6496
rect 5912 6560 6232 6561
rect 5912 6496 5920 6560
rect 5984 6496 6000 6560
rect 6064 6496 6080 6560
rect 6144 6496 6160 6560
rect 6224 6496 6232 6560
rect 5912 6495 6232 6496
rect 2186 6016 2506 6017
rect 2186 5952 2194 6016
rect 2258 5952 2274 6016
rect 2338 5952 2354 6016
rect 2418 5952 2434 6016
rect 2498 5952 2506 6016
rect 2186 5951 2506 5952
rect 4670 6016 4990 6017
rect 4670 5952 4678 6016
rect 4742 5952 4758 6016
rect 4822 5952 4838 6016
rect 4902 5952 4918 6016
rect 4982 5952 4990 6016
rect 4670 5951 4990 5952
rect 7154 6016 7474 6017
rect 7154 5952 7162 6016
rect 7226 5952 7242 6016
rect 7306 5952 7322 6016
rect 7386 5952 7402 6016
rect 7466 5952 7474 6016
rect 7154 5951 7474 5952
rect 7833 5810 7899 5813
rect 8935 5810 9735 5840
rect 7833 5808 9735 5810
rect 7833 5752 7838 5808
rect 7894 5752 9735 5808
rect 7833 5750 9735 5752
rect 7833 5747 7899 5750
rect 8935 5720 9735 5750
rect 3428 5472 3748 5473
rect 3428 5408 3436 5472
rect 3500 5408 3516 5472
rect 3580 5408 3596 5472
rect 3660 5408 3676 5472
rect 3740 5408 3748 5472
rect 3428 5407 3748 5408
rect 5912 5472 6232 5473
rect 5912 5408 5920 5472
rect 5984 5408 6000 5472
rect 6064 5408 6080 5472
rect 6144 5408 6160 5472
rect 6224 5408 6232 5472
rect 5912 5407 6232 5408
rect 2186 4928 2506 4929
rect 2186 4864 2194 4928
rect 2258 4864 2274 4928
rect 2338 4864 2354 4928
rect 2418 4864 2434 4928
rect 2498 4864 2506 4928
rect 2186 4863 2506 4864
rect 4670 4928 4990 4929
rect 4670 4864 4678 4928
rect 4742 4864 4758 4928
rect 4822 4864 4838 4928
rect 4902 4864 4918 4928
rect 4982 4864 4990 4928
rect 4670 4863 4990 4864
rect 7154 4928 7474 4929
rect 7154 4864 7162 4928
rect 7226 4864 7242 4928
rect 7306 4864 7322 4928
rect 7386 4864 7402 4928
rect 7466 4864 7474 4928
rect 7154 4863 7474 4864
rect 3428 4384 3748 4385
rect 3428 4320 3436 4384
rect 3500 4320 3516 4384
rect 3580 4320 3596 4384
rect 3660 4320 3676 4384
rect 3740 4320 3748 4384
rect 3428 4319 3748 4320
rect 5912 4384 6232 4385
rect 5912 4320 5920 4384
rect 5984 4320 6000 4384
rect 6064 4320 6080 4384
rect 6144 4320 6160 4384
rect 6224 4320 6232 4384
rect 5912 4319 6232 4320
rect 0 3906 800 3936
rect 1761 3906 1827 3909
rect 0 3904 1827 3906
rect 0 3848 1766 3904
rect 1822 3848 1827 3904
rect 0 3846 1827 3848
rect 0 3816 800 3846
rect 1761 3843 1827 3846
rect 2186 3840 2506 3841
rect 2186 3776 2194 3840
rect 2258 3776 2274 3840
rect 2338 3776 2354 3840
rect 2418 3776 2434 3840
rect 2498 3776 2506 3840
rect 2186 3775 2506 3776
rect 4670 3840 4990 3841
rect 4670 3776 4678 3840
rect 4742 3776 4758 3840
rect 4822 3776 4838 3840
rect 4902 3776 4918 3840
rect 4982 3776 4990 3840
rect 4670 3775 4990 3776
rect 7154 3840 7474 3841
rect 7154 3776 7162 3840
rect 7226 3776 7242 3840
rect 7306 3776 7322 3840
rect 7386 3776 7402 3840
rect 7466 3776 7474 3840
rect 7154 3775 7474 3776
rect 3428 3296 3748 3297
rect 3428 3232 3436 3296
rect 3500 3232 3516 3296
rect 3580 3232 3596 3296
rect 3660 3232 3676 3296
rect 3740 3232 3748 3296
rect 3428 3231 3748 3232
rect 5912 3296 6232 3297
rect 5912 3232 5920 3296
rect 5984 3232 6000 3296
rect 6064 3232 6080 3296
rect 6144 3232 6160 3296
rect 6224 3232 6232 3296
rect 5912 3231 6232 3232
rect 2186 2752 2506 2753
rect 2186 2688 2194 2752
rect 2258 2688 2274 2752
rect 2338 2688 2354 2752
rect 2418 2688 2434 2752
rect 2498 2688 2506 2752
rect 2186 2687 2506 2688
rect 4670 2752 4990 2753
rect 4670 2688 4678 2752
rect 4742 2688 4758 2752
rect 4822 2688 4838 2752
rect 4902 2688 4918 2752
rect 4982 2688 4990 2752
rect 4670 2687 4990 2688
rect 7154 2752 7474 2753
rect 7154 2688 7162 2752
rect 7226 2688 7242 2752
rect 7306 2688 7322 2752
rect 7386 2688 7402 2752
rect 7466 2688 7474 2752
rect 7154 2687 7474 2688
rect 3428 2208 3748 2209
rect 3428 2144 3436 2208
rect 3500 2144 3516 2208
rect 3580 2144 3596 2208
rect 3660 2144 3676 2208
rect 3740 2144 3748 2208
rect 3428 2143 3748 2144
rect 5912 2208 6232 2209
rect 5912 2144 5920 2208
rect 5984 2144 6000 2208
rect 6064 2144 6080 2208
rect 6144 2144 6160 2208
rect 6224 2144 6232 2208
rect 5912 2143 6232 2144
rect 7741 1730 7807 1733
rect 8935 1730 9735 1760
rect 7741 1728 9735 1730
rect 7741 1672 7746 1728
rect 7802 1672 9735 1728
rect 7741 1670 9735 1672
rect 7741 1667 7807 1670
rect 8935 1640 9735 1670
<< via3 >>
rect 2194 9276 2258 9280
rect 2194 9220 2198 9276
rect 2198 9220 2254 9276
rect 2254 9220 2258 9276
rect 2194 9216 2258 9220
rect 2274 9276 2338 9280
rect 2274 9220 2278 9276
rect 2278 9220 2334 9276
rect 2334 9220 2338 9276
rect 2274 9216 2338 9220
rect 2354 9276 2418 9280
rect 2354 9220 2358 9276
rect 2358 9220 2414 9276
rect 2414 9220 2418 9276
rect 2354 9216 2418 9220
rect 2434 9276 2498 9280
rect 2434 9220 2438 9276
rect 2438 9220 2494 9276
rect 2494 9220 2498 9276
rect 2434 9216 2498 9220
rect 4678 9276 4742 9280
rect 4678 9220 4682 9276
rect 4682 9220 4738 9276
rect 4738 9220 4742 9276
rect 4678 9216 4742 9220
rect 4758 9276 4822 9280
rect 4758 9220 4762 9276
rect 4762 9220 4818 9276
rect 4818 9220 4822 9276
rect 4758 9216 4822 9220
rect 4838 9276 4902 9280
rect 4838 9220 4842 9276
rect 4842 9220 4898 9276
rect 4898 9220 4902 9276
rect 4838 9216 4902 9220
rect 4918 9276 4982 9280
rect 4918 9220 4922 9276
rect 4922 9220 4978 9276
rect 4978 9220 4982 9276
rect 4918 9216 4982 9220
rect 7162 9276 7226 9280
rect 7162 9220 7166 9276
rect 7166 9220 7222 9276
rect 7222 9220 7226 9276
rect 7162 9216 7226 9220
rect 7242 9276 7306 9280
rect 7242 9220 7246 9276
rect 7246 9220 7302 9276
rect 7302 9220 7306 9276
rect 7242 9216 7306 9220
rect 7322 9276 7386 9280
rect 7322 9220 7326 9276
rect 7326 9220 7382 9276
rect 7382 9220 7386 9276
rect 7322 9216 7386 9220
rect 7402 9276 7466 9280
rect 7402 9220 7406 9276
rect 7406 9220 7462 9276
rect 7462 9220 7466 9276
rect 7402 9216 7466 9220
rect 3436 8732 3500 8736
rect 3436 8676 3440 8732
rect 3440 8676 3496 8732
rect 3496 8676 3500 8732
rect 3436 8672 3500 8676
rect 3516 8732 3580 8736
rect 3516 8676 3520 8732
rect 3520 8676 3576 8732
rect 3576 8676 3580 8732
rect 3516 8672 3580 8676
rect 3596 8732 3660 8736
rect 3596 8676 3600 8732
rect 3600 8676 3656 8732
rect 3656 8676 3660 8732
rect 3596 8672 3660 8676
rect 3676 8732 3740 8736
rect 3676 8676 3680 8732
rect 3680 8676 3736 8732
rect 3736 8676 3740 8732
rect 3676 8672 3740 8676
rect 5920 8732 5984 8736
rect 5920 8676 5924 8732
rect 5924 8676 5980 8732
rect 5980 8676 5984 8732
rect 5920 8672 5984 8676
rect 6000 8732 6064 8736
rect 6000 8676 6004 8732
rect 6004 8676 6060 8732
rect 6060 8676 6064 8732
rect 6000 8672 6064 8676
rect 6080 8732 6144 8736
rect 6080 8676 6084 8732
rect 6084 8676 6140 8732
rect 6140 8676 6144 8732
rect 6080 8672 6144 8676
rect 6160 8732 6224 8736
rect 6160 8676 6164 8732
rect 6164 8676 6220 8732
rect 6220 8676 6224 8732
rect 6160 8672 6224 8676
rect 2194 8188 2258 8192
rect 2194 8132 2198 8188
rect 2198 8132 2254 8188
rect 2254 8132 2258 8188
rect 2194 8128 2258 8132
rect 2274 8188 2338 8192
rect 2274 8132 2278 8188
rect 2278 8132 2334 8188
rect 2334 8132 2338 8188
rect 2274 8128 2338 8132
rect 2354 8188 2418 8192
rect 2354 8132 2358 8188
rect 2358 8132 2414 8188
rect 2414 8132 2418 8188
rect 2354 8128 2418 8132
rect 2434 8188 2498 8192
rect 2434 8132 2438 8188
rect 2438 8132 2494 8188
rect 2494 8132 2498 8188
rect 2434 8128 2498 8132
rect 4678 8188 4742 8192
rect 4678 8132 4682 8188
rect 4682 8132 4738 8188
rect 4738 8132 4742 8188
rect 4678 8128 4742 8132
rect 4758 8188 4822 8192
rect 4758 8132 4762 8188
rect 4762 8132 4818 8188
rect 4818 8132 4822 8188
rect 4758 8128 4822 8132
rect 4838 8188 4902 8192
rect 4838 8132 4842 8188
rect 4842 8132 4898 8188
rect 4898 8132 4902 8188
rect 4838 8128 4902 8132
rect 4918 8188 4982 8192
rect 4918 8132 4922 8188
rect 4922 8132 4978 8188
rect 4978 8132 4982 8188
rect 4918 8128 4982 8132
rect 7162 8188 7226 8192
rect 7162 8132 7166 8188
rect 7166 8132 7222 8188
rect 7222 8132 7226 8188
rect 7162 8128 7226 8132
rect 7242 8188 7306 8192
rect 7242 8132 7246 8188
rect 7246 8132 7302 8188
rect 7302 8132 7306 8188
rect 7242 8128 7306 8132
rect 7322 8188 7386 8192
rect 7322 8132 7326 8188
rect 7326 8132 7382 8188
rect 7382 8132 7386 8188
rect 7322 8128 7386 8132
rect 7402 8188 7466 8192
rect 7402 8132 7406 8188
rect 7406 8132 7462 8188
rect 7462 8132 7466 8188
rect 7402 8128 7466 8132
rect 3436 7644 3500 7648
rect 3436 7588 3440 7644
rect 3440 7588 3496 7644
rect 3496 7588 3500 7644
rect 3436 7584 3500 7588
rect 3516 7644 3580 7648
rect 3516 7588 3520 7644
rect 3520 7588 3576 7644
rect 3576 7588 3580 7644
rect 3516 7584 3580 7588
rect 3596 7644 3660 7648
rect 3596 7588 3600 7644
rect 3600 7588 3656 7644
rect 3656 7588 3660 7644
rect 3596 7584 3660 7588
rect 3676 7644 3740 7648
rect 3676 7588 3680 7644
rect 3680 7588 3736 7644
rect 3736 7588 3740 7644
rect 3676 7584 3740 7588
rect 5920 7644 5984 7648
rect 5920 7588 5924 7644
rect 5924 7588 5980 7644
rect 5980 7588 5984 7644
rect 5920 7584 5984 7588
rect 6000 7644 6064 7648
rect 6000 7588 6004 7644
rect 6004 7588 6060 7644
rect 6060 7588 6064 7644
rect 6000 7584 6064 7588
rect 6080 7644 6144 7648
rect 6080 7588 6084 7644
rect 6084 7588 6140 7644
rect 6140 7588 6144 7644
rect 6080 7584 6144 7588
rect 6160 7644 6224 7648
rect 6160 7588 6164 7644
rect 6164 7588 6220 7644
rect 6220 7588 6224 7644
rect 6160 7584 6224 7588
rect 2194 7100 2258 7104
rect 2194 7044 2198 7100
rect 2198 7044 2254 7100
rect 2254 7044 2258 7100
rect 2194 7040 2258 7044
rect 2274 7100 2338 7104
rect 2274 7044 2278 7100
rect 2278 7044 2334 7100
rect 2334 7044 2338 7100
rect 2274 7040 2338 7044
rect 2354 7100 2418 7104
rect 2354 7044 2358 7100
rect 2358 7044 2414 7100
rect 2414 7044 2418 7100
rect 2354 7040 2418 7044
rect 2434 7100 2498 7104
rect 2434 7044 2438 7100
rect 2438 7044 2494 7100
rect 2494 7044 2498 7100
rect 2434 7040 2498 7044
rect 4678 7100 4742 7104
rect 4678 7044 4682 7100
rect 4682 7044 4738 7100
rect 4738 7044 4742 7100
rect 4678 7040 4742 7044
rect 4758 7100 4822 7104
rect 4758 7044 4762 7100
rect 4762 7044 4818 7100
rect 4818 7044 4822 7100
rect 4758 7040 4822 7044
rect 4838 7100 4902 7104
rect 4838 7044 4842 7100
rect 4842 7044 4898 7100
rect 4898 7044 4902 7100
rect 4838 7040 4902 7044
rect 4918 7100 4982 7104
rect 4918 7044 4922 7100
rect 4922 7044 4978 7100
rect 4978 7044 4982 7100
rect 4918 7040 4982 7044
rect 7162 7100 7226 7104
rect 7162 7044 7166 7100
rect 7166 7044 7222 7100
rect 7222 7044 7226 7100
rect 7162 7040 7226 7044
rect 7242 7100 7306 7104
rect 7242 7044 7246 7100
rect 7246 7044 7302 7100
rect 7302 7044 7306 7100
rect 7242 7040 7306 7044
rect 7322 7100 7386 7104
rect 7322 7044 7326 7100
rect 7326 7044 7382 7100
rect 7382 7044 7386 7100
rect 7322 7040 7386 7044
rect 7402 7100 7466 7104
rect 7402 7044 7406 7100
rect 7406 7044 7462 7100
rect 7462 7044 7466 7100
rect 7402 7040 7466 7044
rect 3436 6556 3500 6560
rect 3436 6500 3440 6556
rect 3440 6500 3496 6556
rect 3496 6500 3500 6556
rect 3436 6496 3500 6500
rect 3516 6556 3580 6560
rect 3516 6500 3520 6556
rect 3520 6500 3576 6556
rect 3576 6500 3580 6556
rect 3516 6496 3580 6500
rect 3596 6556 3660 6560
rect 3596 6500 3600 6556
rect 3600 6500 3656 6556
rect 3656 6500 3660 6556
rect 3596 6496 3660 6500
rect 3676 6556 3740 6560
rect 3676 6500 3680 6556
rect 3680 6500 3736 6556
rect 3736 6500 3740 6556
rect 3676 6496 3740 6500
rect 5920 6556 5984 6560
rect 5920 6500 5924 6556
rect 5924 6500 5980 6556
rect 5980 6500 5984 6556
rect 5920 6496 5984 6500
rect 6000 6556 6064 6560
rect 6000 6500 6004 6556
rect 6004 6500 6060 6556
rect 6060 6500 6064 6556
rect 6000 6496 6064 6500
rect 6080 6556 6144 6560
rect 6080 6500 6084 6556
rect 6084 6500 6140 6556
rect 6140 6500 6144 6556
rect 6080 6496 6144 6500
rect 6160 6556 6224 6560
rect 6160 6500 6164 6556
rect 6164 6500 6220 6556
rect 6220 6500 6224 6556
rect 6160 6496 6224 6500
rect 2194 6012 2258 6016
rect 2194 5956 2198 6012
rect 2198 5956 2254 6012
rect 2254 5956 2258 6012
rect 2194 5952 2258 5956
rect 2274 6012 2338 6016
rect 2274 5956 2278 6012
rect 2278 5956 2334 6012
rect 2334 5956 2338 6012
rect 2274 5952 2338 5956
rect 2354 6012 2418 6016
rect 2354 5956 2358 6012
rect 2358 5956 2414 6012
rect 2414 5956 2418 6012
rect 2354 5952 2418 5956
rect 2434 6012 2498 6016
rect 2434 5956 2438 6012
rect 2438 5956 2494 6012
rect 2494 5956 2498 6012
rect 2434 5952 2498 5956
rect 4678 6012 4742 6016
rect 4678 5956 4682 6012
rect 4682 5956 4738 6012
rect 4738 5956 4742 6012
rect 4678 5952 4742 5956
rect 4758 6012 4822 6016
rect 4758 5956 4762 6012
rect 4762 5956 4818 6012
rect 4818 5956 4822 6012
rect 4758 5952 4822 5956
rect 4838 6012 4902 6016
rect 4838 5956 4842 6012
rect 4842 5956 4898 6012
rect 4898 5956 4902 6012
rect 4838 5952 4902 5956
rect 4918 6012 4982 6016
rect 4918 5956 4922 6012
rect 4922 5956 4978 6012
rect 4978 5956 4982 6012
rect 4918 5952 4982 5956
rect 7162 6012 7226 6016
rect 7162 5956 7166 6012
rect 7166 5956 7222 6012
rect 7222 5956 7226 6012
rect 7162 5952 7226 5956
rect 7242 6012 7306 6016
rect 7242 5956 7246 6012
rect 7246 5956 7302 6012
rect 7302 5956 7306 6012
rect 7242 5952 7306 5956
rect 7322 6012 7386 6016
rect 7322 5956 7326 6012
rect 7326 5956 7382 6012
rect 7382 5956 7386 6012
rect 7322 5952 7386 5956
rect 7402 6012 7466 6016
rect 7402 5956 7406 6012
rect 7406 5956 7462 6012
rect 7462 5956 7466 6012
rect 7402 5952 7466 5956
rect 3436 5468 3500 5472
rect 3436 5412 3440 5468
rect 3440 5412 3496 5468
rect 3496 5412 3500 5468
rect 3436 5408 3500 5412
rect 3516 5468 3580 5472
rect 3516 5412 3520 5468
rect 3520 5412 3576 5468
rect 3576 5412 3580 5468
rect 3516 5408 3580 5412
rect 3596 5468 3660 5472
rect 3596 5412 3600 5468
rect 3600 5412 3656 5468
rect 3656 5412 3660 5468
rect 3596 5408 3660 5412
rect 3676 5468 3740 5472
rect 3676 5412 3680 5468
rect 3680 5412 3736 5468
rect 3736 5412 3740 5468
rect 3676 5408 3740 5412
rect 5920 5468 5984 5472
rect 5920 5412 5924 5468
rect 5924 5412 5980 5468
rect 5980 5412 5984 5468
rect 5920 5408 5984 5412
rect 6000 5468 6064 5472
rect 6000 5412 6004 5468
rect 6004 5412 6060 5468
rect 6060 5412 6064 5468
rect 6000 5408 6064 5412
rect 6080 5468 6144 5472
rect 6080 5412 6084 5468
rect 6084 5412 6140 5468
rect 6140 5412 6144 5468
rect 6080 5408 6144 5412
rect 6160 5468 6224 5472
rect 6160 5412 6164 5468
rect 6164 5412 6220 5468
rect 6220 5412 6224 5468
rect 6160 5408 6224 5412
rect 2194 4924 2258 4928
rect 2194 4868 2198 4924
rect 2198 4868 2254 4924
rect 2254 4868 2258 4924
rect 2194 4864 2258 4868
rect 2274 4924 2338 4928
rect 2274 4868 2278 4924
rect 2278 4868 2334 4924
rect 2334 4868 2338 4924
rect 2274 4864 2338 4868
rect 2354 4924 2418 4928
rect 2354 4868 2358 4924
rect 2358 4868 2414 4924
rect 2414 4868 2418 4924
rect 2354 4864 2418 4868
rect 2434 4924 2498 4928
rect 2434 4868 2438 4924
rect 2438 4868 2494 4924
rect 2494 4868 2498 4924
rect 2434 4864 2498 4868
rect 4678 4924 4742 4928
rect 4678 4868 4682 4924
rect 4682 4868 4738 4924
rect 4738 4868 4742 4924
rect 4678 4864 4742 4868
rect 4758 4924 4822 4928
rect 4758 4868 4762 4924
rect 4762 4868 4818 4924
rect 4818 4868 4822 4924
rect 4758 4864 4822 4868
rect 4838 4924 4902 4928
rect 4838 4868 4842 4924
rect 4842 4868 4898 4924
rect 4898 4868 4902 4924
rect 4838 4864 4902 4868
rect 4918 4924 4982 4928
rect 4918 4868 4922 4924
rect 4922 4868 4978 4924
rect 4978 4868 4982 4924
rect 4918 4864 4982 4868
rect 7162 4924 7226 4928
rect 7162 4868 7166 4924
rect 7166 4868 7222 4924
rect 7222 4868 7226 4924
rect 7162 4864 7226 4868
rect 7242 4924 7306 4928
rect 7242 4868 7246 4924
rect 7246 4868 7302 4924
rect 7302 4868 7306 4924
rect 7242 4864 7306 4868
rect 7322 4924 7386 4928
rect 7322 4868 7326 4924
rect 7326 4868 7382 4924
rect 7382 4868 7386 4924
rect 7322 4864 7386 4868
rect 7402 4924 7466 4928
rect 7402 4868 7406 4924
rect 7406 4868 7462 4924
rect 7462 4868 7466 4924
rect 7402 4864 7466 4868
rect 3436 4380 3500 4384
rect 3436 4324 3440 4380
rect 3440 4324 3496 4380
rect 3496 4324 3500 4380
rect 3436 4320 3500 4324
rect 3516 4380 3580 4384
rect 3516 4324 3520 4380
rect 3520 4324 3576 4380
rect 3576 4324 3580 4380
rect 3516 4320 3580 4324
rect 3596 4380 3660 4384
rect 3596 4324 3600 4380
rect 3600 4324 3656 4380
rect 3656 4324 3660 4380
rect 3596 4320 3660 4324
rect 3676 4380 3740 4384
rect 3676 4324 3680 4380
rect 3680 4324 3736 4380
rect 3736 4324 3740 4380
rect 3676 4320 3740 4324
rect 5920 4380 5984 4384
rect 5920 4324 5924 4380
rect 5924 4324 5980 4380
rect 5980 4324 5984 4380
rect 5920 4320 5984 4324
rect 6000 4380 6064 4384
rect 6000 4324 6004 4380
rect 6004 4324 6060 4380
rect 6060 4324 6064 4380
rect 6000 4320 6064 4324
rect 6080 4380 6144 4384
rect 6080 4324 6084 4380
rect 6084 4324 6140 4380
rect 6140 4324 6144 4380
rect 6080 4320 6144 4324
rect 6160 4380 6224 4384
rect 6160 4324 6164 4380
rect 6164 4324 6220 4380
rect 6220 4324 6224 4380
rect 6160 4320 6224 4324
rect 2194 3836 2258 3840
rect 2194 3780 2198 3836
rect 2198 3780 2254 3836
rect 2254 3780 2258 3836
rect 2194 3776 2258 3780
rect 2274 3836 2338 3840
rect 2274 3780 2278 3836
rect 2278 3780 2334 3836
rect 2334 3780 2338 3836
rect 2274 3776 2338 3780
rect 2354 3836 2418 3840
rect 2354 3780 2358 3836
rect 2358 3780 2414 3836
rect 2414 3780 2418 3836
rect 2354 3776 2418 3780
rect 2434 3836 2498 3840
rect 2434 3780 2438 3836
rect 2438 3780 2494 3836
rect 2494 3780 2498 3836
rect 2434 3776 2498 3780
rect 4678 3836 4742 3840
rect 4678 3780 4682 3836
rect 4682 3780 4738 3836
rect 4738 3780 4742 3836
rect 4678 3776 4742 3780
rect 4758 3836 4822 3840
rect 4758 3780 4762 3836
rect 4762 3780 4818 3836
rect 4818 3780 4822 3836
rect 4758 3776 4822 3780
rect 4838 3836 4902 3840
rect 4838 3780 4842 3836
rect 4842 3780 4898 3836
rect 4898 3780 4902 3836
rect 4838 3776 4902 3780
rect 4918 3836 4982 3840
rect 4918 3780 4922 3836
rect 4922 3780 4978 3836
rect 4978 3780 4982 3836
rect 4918 3776 4982 3780
rect 7162 3836 7226 3840
rect 7162 3780 7166 3836
rect 7166 3780 7222 3836
rect 7222 3780 7226 3836
rect 7162 3776 7226 3780
rect 7242 3836 7306 3840
rect 7242 3780 7246 3836
rect 7246 3780 7302 3836
rect 7302 3780 7306 3836
rect 7242 3776 7306 3780
rect 7322 3836 7386 3840
rect 7322 3780 7326 3836
rect 7326 3780 7382 3836
rect 7382 3780 7386 3836
rect 7322 3776 7386 3780
rect 7402 3836 7466 3840
rect 7402 3780 7406 3836
rect 7406 3780 7462 3836
rect 7462 3780 7466 3836
rect 7402 3776 7466 3780
rect 3436 3292 3500 3296
rect 3436 3236 3440 3292
rect 3440 3236 3496 3292
rect 3496 3236 3500 3292
rect 3436 3232 3500 3236
rect 3516 3292 3580 3296
rect 3516 3236 3520 3292
rect 3520 3236 3576 3292
rect 3576 3236 3580 3292
rect 3516 3232 3580 3236
rect 3596 3292 3660 3296
rect 3596 3236 3600 3292
rect 3600 3236 3656 3292
rect 3656 3236 3660 3292
rect 3596 3232 3660 3236
rect 3676 3292 3740 3296
rect 3676 3236 3680 3292
rect 3680 3236 3736 3292
rect 3736 3236 3740 3292
rect 3676 3232 3740 3236
rect 5920 3292 5984 3296
rect 5920 3236 5924 3292
rect 5924 3236 5980 3292
rect 5980 3236 5984 3292
rect 5920 3232 5984 3236
rect 6000 3292 6064 3296
rect 6000 3236 6004 3292
rect 6004 3236 6060 3292
rect 6060 3236 6064 3292
rect 6000 3232 6064 3236
rect 6080 3292 6144 3296
rect 6080 3236 6084 3292
rect 6084 3236 6140 3292
rect 6140 3236 6144 3292
rect 6080 3232 6144 3236
rect 6160 3292 6224 3296
rect 6160 3236 6164 3292
rect 6164 3236 6220 3292
rect 6220 3236 6224 3292
rect 6160 3232 6224 3236
rect 2194 2748 2258 2752
rect 2194 2692 2198 2748
rect 2198 2692 2254 2748
rect 2254 2692 2258 2748
rect 2194 2688 2258 2692
rect 2274 2748 2338 2752
rect 2274 2692 2278 2748
rect 2278 2692 2334 2748
rect 2334 2692 2338 2748
rect 2274 2688 2338 2692
rect 2354 2748 2418 2752
rect 2354 2692 2358 2748
rect 2358 2692 2414 2748
rect 2414 2692 2418 2748
rect 2354 2688 2418 2692
rect 2434 2748 2498 2752
rect 2434 2692 2438 2748
rect 2438 2692 2494 2748
rect 2494 2692 2498 2748
rect 2434 2688 2498 2692
rect 4678 2748 4742 2752
rect 4678 2692 4682 2748
rect 4682 2692 4738 2748
rect 4738 2692 4742 2748
rect 4678 2688 4742 2692
rect 4758 2748 4822 2752
rect 4758 2692 4762 2748
rect 4762 2692 4818 2748
rect 4818 2692 4822 2748
rect 4758 2688 4822 2692
rect 4838 2748 4902 2752
rect 4838 2692 4842 2748
rect 4842 2692 4898 2748
rect 4898 2692 4902 2748
rect 4838 2688 4902 2692
rect 4918 2748 4982 2752
rect 4918 2692 4922 2748
rect 4922 2692 4978 2748
rect 4978 2692 4982 2748
rect 4918 2688 4982 2692
rect 7162 2748 7226 2752
rect 7162 2692 7166 2748
rect 7166 2692 7222 2748
rect 7222 2692 7226 2748
rect 7162 2688 7226 2692
rect 7242 2748 7306 2752
rect 7242 2692 7246 2748
rect 7246 2692 7302 2748
rect 7302 2692 7306 2748
rect 7242 2688 7306 2692
rect 7322 2748 7386 2752
rect 7322 2692 7326 2748
rect 7326 2692 7382 2748
rect 7382 2692 7386 2748
rect 7322 2688 7386 2692
rect 7402 2748 7466 2752
rect 7402 2692 7406 2748
rect 7406 2692 7462 2748
rect 7462 2692 7466 2748
rect 7402 2688 7466 2692
rect 3436 2204 3500 2208
rect 3436 2148 3440 2204
rect 3440 2148 3496 2204
rect 3496 2148 3500 2204
rect 3436 2144 3500 2148
rect 3516 2204 3580 2208
rect 3516 2148 3520 2204
rect 3520 2148 3576 2204
rect 3576 2148 3580 2204
rect 3516 2144 3580 2148
rect 3596 2204 3660 2208
rect 3596 2148 3600 2204
rect 3600 2148 3656 2204
rect 3656 2148 3660 2204
rect 3596 2144 3660 2148
rect 3676 2204 3740 2208
rect 3676 2148 3680 2204
rect 3680 2148 3736 2204
rect 3736 2148 3740 2204
rect 3676 2144 3740 2148
rect 5920 2204 5984 2208
rect 5920 2148 5924 2204
rect 5924 2148 5980 2204
rect 5980 2148 5984 2204
rect 5920 2144 5984 2148
rect 6000 2204 6064 2208
rect 6000 2148 6004 2204
rect 6004 2148 6060 2204
rect 6060 2148 6064 2204
rect 6000 2144 6064 2148
rect 6080 2204 6144 2208
rect 6080 2148 6084 2204
rect 6084 2148 6140 2204
rect 6140 2148 6144 2204
rect 6080 2144 6144 2148
rect 6160 2204 6224 2208
rect 6160 2148 6164 2204
rect 6164 2148 6220 2204
rect 6220 2148 6224 2204
rect 6160 2144 6224 2148
<< metal4 >>
rect 2186 9280 2506 9296
rect 2186 9216 2194 9280
rect 2258 9216 2274 9280
rect 2338 9216 2354 9280
rect 2418 9216 2434 9280
rect 2498 9216 2506 9280
rect 2186 8192 2506 9216
rect 2186 8128 2194 8192
rect 2258 8139 2274 8192
rect 2338 8139 2354 8192
rect 2418 8139 2434 8192
rect 2498 8128 2506 8192
rect 2186 7903 2228 8128
rect 2464 7903 2506 8128
rect 2186 7104 2506 7903
rect 2186 7040 2194 7104
rect 2258 7040 2274 7104
rect 2338 7040 2354 7104
rect 2418 7040 2434 7104
rect 2498 7040 2506 7104
rect 2186 6016 2506 7040
rect 2186 5952 2194 6016
rect 2258 5952 2274 6016
rect 2338 5952 2354 6016
rect 2418 5952 2434 6016
rect 2498 5952 2506 6016
rect 2186 5782 2506 5952
rect 2186 5546 2228 5782
rect 2464 5546 2506 5782
rect 2186 4928 2506 5546
rect 2186 4864 2194 4928
rect 2258 4864 2274 4928
rect 2338 4864 2354 4928
rect 2418 4864 2434 4928
rect 2498 4864 2506 4928
rect 2186 3840 2506 4864
rect 2186 3776 2194 3840
rect 2258 3776 2274 3840
rect 2338 3776 2354 3840
rect 2418 3776 2434 3840
rect 2498 3776 2506 3840
rect 2186 3424 2506 3776
rect 2186 3188 2228 3424
rect 2464 3188 2506 3424
rect 2186 2752 2506 3188
rect 2186 2688 2194 2752
rect 2258 2688 2274 2752
rect 2338 2688 2354 2752
rect 2418 2688 2434 2752
rect 2498 2688 2506 2752
rect 2186 2128 2506 2688
rect 3428 8736 3748 9296
rect 3428 8672 3436 8736
rect 3500 8672 3516 8736
rect 3580 8672 3596 8736
rect 3660 8672 3676 8736
rect 3740 8672 3748 8736
rect 3428 7648 3748 8672
rect 3428 7584 3436 7648
rect 3500 7584 3516 7648
rect 3580 7584 3596 7648
rect 3660 7584 3676 7648
rect 3740 7584 3748 7648
rect 3428 6960 3748 7584
rect 3428 6724 3470 6960
rect 3706 6724 3748 6960
rect 3428 6560 3748 6724
rect 3428 6496 3436 6560
rect 3500 6496 3516 6560
rect 3580 6496 3596 6560
rect 3660 6496 3676 6560
rect 3740 6496 3748 6560
rect 3428 5472 3748 6496
rect 3428 5408 3436 5472
rect 3500 5408 3516 5472
rect 3580 5408 3596 5472
rect 3660 5408 3676 5472
rect 3740 5408 3748 5472
rect 3428 4603 3748 5408
rect 3428 4384 3470 4603
rect 3706 4384 3748 4603
rect 3428 4320 3436 4384
rect 3500 4320 3516 4367
rect 3580 4320 3596 4367
rect 3660 4320 3676 4367
rect 3740 4320 3748 4384
rect 3428 3296 3748 4320
rect 3428 3232 3436 3296
rect 3500 3232 3516 3296
rect 3580 3232 3596 3296
rect 3660 3232 3676 3296
rect 3740 3232 3748 3296
rect 3428 2208 3748 3232
rect 3428 2144 3436 2208
rect 3500 2144 3516 2208
rect 3580 2144 3596 2208
rect 3660 2144 3676 2208
rect 3740 2144 3748 2208
rect 3428 2128 3748 2144
rect 4670 9280 4990 9296
rect 4670 9216 4678 9280
rect 4742 9216 4758 9280
rect 4822 9216 4838 9280
rect 4902 9216 4918 9280
rect 4982 9216 4990 9280
rect 4670 8192 4990 9216
rect 4670 8128 4678 8192
rect 4742 8139 4758 8192
rect 4822 8139 4838 8192
rect 4902 8139 4918 8192
rect 4982 8128 4990 8192
rect 4670 7903 4712 8128
rect 4948 7903 4990 8128
rect 4670 7104 4990 7903
rect 4670 7040 4678 7104
rect 4742 7040 4758 7104
rect 4822 7040 4838 7104
rect 4902 7040 4918 7104
rect 4982 7040 4990 7104
rect 4670 6016 4990 7040
rect 4670 5952 4678 6016
rect 4742 5952 4758 6016
rect 4822 5952 4838 6016
rect 4902 5952 4918 6016
rect 4982 5952 4990 6016
rect 4670 5782 4990 5952
rect 4670 5546 4712 5782
rect 4948 5546 4990 5782
rect 4670 4928 4990 5546
rect 4670 4864 4678 4928
rect 4742 4864 4758 4928
rect 4822 4864 4838 4928
rect 4902 4864 4918 4928
rect 4982 4864 4990 4928
rect 4670 3840 4990 4864
rect 4670 3776 4678 3840
rect 4742 3776 4758 3840
rect 4822 3776 4838 3840
rect 4902 3776 4918 3840
rect 4982 3776 4990 3840
rect 4670 3424 4990 3776
rect 4670 3188 4712 3424
rect 4948 3188 4990 3424
rect 4670 2752 4990 3188
rect 4670 2688 4678 2752
rect 4742 2688 4758 2752
rect 4822 2688 4838 2752
rect 4902 2688 4918 2752
rect 4982 2688 4990 2752
rect 4670 2128 4990 2688
rect 5912 8736 6232 9296
rect 5912 8672 5920 8736
rect 5984 8672 6000 8736
rect 6064 8672 6080 8736
rect 6144 8672 6160 8736
rect 6224 8672 6232 8736
rect 5912 7648 6232 8672
rect 5912 7584 5920 7648
rect 5984 7584 6000 7648
rect 6064 7584 6080 7648
rect 6144 7584 6160 7648
rect 6224 7584 6232 7648
rect 5912 6960 6232 7584
rect 5912 6724 5954 6960
rect 6190 6724 6232 6960
rect 5912 6560 6232 6724
rect 5912 6496 5920 6560
rect 5984 6496 6000 6560
rect 6064 6496 6080 6560
rect 6144 6496 6160 6560
rect 6224 6496 6232 6560
rect 5912 5472 6232 6496
rect 5912 5408 5920 5472
rect 5984 5408 6000 5472
rect 6064 5408 6080 5472
rect 6144 5408 6160 5472
rect 6224 5408 6232 5472
rect 5912 4603 6232 5408
rect 5912 4384 5954 4603
rect 6190 4384 6232 4603
rect 5912 4320 5920 4384
rect 5984 4320 6000 4367
rect 6064 4320 6080 4367
rect 6144 4320 6160 4367
rect 6224 4320 6232 4384
rect 5912 3296 6232 4320
rect 5912 3232 5920 3296
rect 5984 3232 6000 3296
rect 6064 3232 6080 3296
rect 6144 3232 6160 3296
rect 6224 3232 6232 3296
rect 5912 2208 6232 3232
rect 5912 2144 5920 2208
rect 5984 2144 6000 2208
rect 6064 2144 6080 2208
rect 6144 2144 6160 2208
rect 6224 2144 6232 2208
rect 5912 2128 6232 2144
rect 7154 9280 7474 9296
rect 7154 9216 7162 9280
rect 7226 9216 7242 9280
rect 7306 9216 7322 9280
rect 7386 9216 7402 9280
rect 7466 9216 7474 9280
rect 7154 8192 7474 9216
rect 7154 8128 7162 8192
rect 7226 8139 7242 8192
rect 7306 8139 7322 8192
rect 7386 8139 7402 8192
rect 7466 8128 7474 8192
rect 7154 7903 7196 8128
rect 7432 7903 7474 8128
rect 7154 7104 7474 7903
rect 7154 7040 7162 7104
rect 7226 7040 7242 7104
rect 7306 7040 7322 7104
rect 7386 7040 7402 7104
rect 7466 7040 7474 7104
rect 7154 6016 7474 7040
rect 7154 5952 7162 6016
rect 7226 5952 7242 6016
rect 7306 5952 7322 6016
rect 7386 5952 7402 6016
rect 7466 5952 7474 6016
rect 7154 5782 7474 5952
rect 7154 5546 7196 5782
rect 7432 5546 7474 5782
rect 7154 4928 7474 5546
rect 7154 4864 7162 4928
rect 7226 4864 7242 4928
rect 7306 4864 7322 4928
rect 7386 4864 7402 4928
rect 7466 4864 7474 4928
rect 7154 3840 7474 4864
rect 7154 3776 7162 3840
rect 7226 3776 7242 3840
rect 7306 3776 7322 3840
rect 7386 3776 7402 3840
rect 7466 3776 7474 3840
rect 7154 3424 7474 3776
rect 7154 3188 7196 3424
rect 7432 3188 7474 3424
rect 7154 2752 7474 3188
rect 7154 2688 7162 2752
rect 7226 2688 7242 2752
rect 7306 2688 7322 2752
rect 7386 2688 7402 2752
rect 7466 2688 7474 2752
rect 7154 2128 7474 2688
<< via4 >>
rect 2228 8128 2258 8139
rect 2258 8128 2274 8139
rect 2274 8128 2338 8139
rect 2338 8128 2354 8139
rect 2354 8128 2418 8139
rect 2418 8128 2434 8139
rect 2434 8128 2464 8139
rect 2228 7903 2464 8128
rect 2228 5546 2464 5782
rect 2228 3188 2464 3424
rect 3470 6724 3706 6960
rect 3470 4384 3706 4603
rect 3470 4367 3500 4384
rect 3500 4367 3516 4384
rect 3516 4367 3580 4384
rect 3580 4367 3596 4384
rect 3596 4367 3660 4384
rect 3660 4367 3676 4384
rect 3676 4367 3706 4384
rect 4712 8128 4742 8139
rect 4742 8128 4758 8139
rect 4758 8128 4822 8139
rect 4822 8128 4838 8139
rect 4838 8128 4902 8139
rect 4902 8128 4918 8139
rect 4918 8128 4948 8139
rect 4712 7903 4948 8128
rect 4712 5546 4948 5782
rect 4712 3188 4948 3424
rect 5954 6724 6190 6960
rect 5954 4384 6190 4603
rect 5954 4367 5984 4384
rect 5984 4367 6000 4384
rect 6000 4367 6064 4384
rect 6064 4367 6080 4384
rect 6080 4367 6144 4384
rect 6144 4367 6160 4384
rect 6160 4367 6190 4384
rect 7196 8128 7226 8139
rect 7226 8128 7242 8139
rect 7242 8128 7306 8139
rect 7306 8128 7322 8139
rect 7322 8128 7386 8139
rect 7386 8128 7402 8139
rect 7402 8128 7432 8139
rect 7196 7903 7432 8128
rect 7196 5546 7432 5782
rect 7196 3188 7432 3424
<< metal5 >>
rect 1104 8139 8556 8181
rect 1104 7903 2228 8139
rect 2464 7903 4712 8139
rect 4948 7903 7196 8139
rect 7432 7903 8556 8139
rect 1104 7861 8556 7903
rect 1104 6960 8556 7002
rect 1104 6724 3470 6960
rect 3706 6724 5954 6960
rect 6190 6724 8556 6960
rect 1104 6682 8556 6724
rect 1104 5782 8556 5824
rect 1104 5546 2228 5782
rect 2464 5546 4712 5782
rect 4948 5546 7196 5782
rect 7432 5546 8556 5782
rect 1104 5504 8556 5546
rect 1104 4603 8556 4646
rect 1104 4367 3470 4603
rect 3706 4367 5954 4603
rect 6190 4367 8556 4603
rect 1104 4325 8556 4367
rect 1104 3424 8556 3466
rect 1104 3188 2228 3424
rect 2464 3188 4712 3424
rect 4948 3188 7196 3424
rect 7432 3188 8556 3424
rect 1104 3146 8556 3188
use sky130_fd_sc_hd__clkbuf_1  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform -1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1629961164
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform 1 0 2024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1629961164
transform -1 0 2944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform 1 0 2576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1629961164
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1629961164
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41
timestamp 1629961164
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1629961164
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1629961164
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50
timestamp 1629961164
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1629961164
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1629961164
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1629961164
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1629961164
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1629961164
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1629961164
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1629961164
transform -1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65
timestamp 1629961164
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1629961164
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform 1 0 7452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1629961164
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1629961164
transform -1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1629961164
transform -1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform -1 0 7912 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1629961164
transform 1 0 7636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1629961164
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1629961164
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1629961164
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1629961164
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1629961164
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1629961164
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1629961164
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1629961164
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1629961164
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_77
timestamp 1629961164
transform 1 0 8188 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1629961164
transform -1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_10
timestamp 1629961164
transform 1 0 2024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1629961164
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1629961164
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1629961164
transform -1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_22
timestamp 1629961164
transform 1 0 3128 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_34
timestamp 1629961164
transform 1 0 4232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_46
timestamp 1629961164
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1629961164
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1629961164
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1629961164
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_69
timestamp 1629961164
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_77
timestamp 1629961164
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1629961164
transform -1 0 8556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1629961164
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1629961164
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1629961164
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1629961164
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1629961164
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_41
timestamp 1629961164
transform 1 0 4876 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1629961164
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_47
timestamp 1629961164
transform 1 0 5428 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_59
timestamp 1629961164
transform 1 0 6532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _12_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform -1 0 5428 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_4_71
timestamp 1629961164
transform 1 0 7636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_77
timestamp 1629961164
transform 1 0 8188 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1629961164
transform -1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1629961164
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1629961164
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1629961164
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _16_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform -1 0 2484 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform 1 0 2852 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_35
timestamp 1629961164
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _17_
timestamp 1629961164
transform 1 0 4692 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1629961164
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1629961164
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1629961164
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_69
timestamp 1629961164
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_77
timestamp 1629961164
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1629961164
transform -1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1629961164
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1629961164
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1629961164
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1629961164
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1629961164
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _15_
timestamp 1629961164
transform 1 0 2852 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform -1 0 3312 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1629961164
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_28
timestamp 1629961164
transform 1 0 3680 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1629961164
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _23_
timestamp 1629961164
transform 1 0 3772 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _32_
timestamp 1629961164
transform 1 0 4416 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_45
timestamp 1629961164
transform 1 0 5244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_58
timestamp 1629961164
transform 1 0 6440 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1629961164
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1629961164
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _13_
timestamp 1629961164
transform -1 0 6440 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _18_
timestamp 1629961164
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_70
timestamp 1629961164
transform 1 0 7544 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_66
timestamp 1629961164
transform 1 0 7176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1629961164
transform 1 0 7544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_74
timestamp 1629961164
transform 1 0 7912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1629961164
transform -1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1629961164
transform -1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1629961164
transform 1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1629961164
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1629961164
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1629961164
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _30_
timestamp 1629961164
transform -1 0 3312 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1629961164
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1629961164
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1629961164
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _24_
timestamp 1629961164
transform 1 0 3864 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_46
timestamp 1629961164
transform 1 0 5336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _28_
timestamp 1629961164
transform 1 0 5704 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1629961164
transform 1 0 7176 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1629961164
transform -1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1629961164
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1629961164
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1629961164
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _29_
timestamp 1629961164
transform 1 0 2024 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_9_26
timestamp 1629961164
transform 1 0 3496 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1629961164
transform 1 0 4048 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1629961164
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1629961164
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _14_
timestamp 1629961164
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_66
timestamp 1629961164
transform 1 0 7176 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1629961164
transform -1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1629961164
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1629961164
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1629961164
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _31_
timestamp 1629961164
transform -1 0 3312 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1629961164
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_38
timestamp 1629961164
transform 1 0 4600 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1629961164
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _21_
timestamp 1629961164
transform 1 0 3772 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_44
timestamp 1629961164
transform 1 0 5152 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1629961164
transform 1 0 5244 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_10_65
timestamp 1629961164
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_74
timestamp 1629961164
transform 1 0 7912 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1629961164
transform -1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1629961164
transform 1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1629961164
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_9
timestamp 1629961164
transform 1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1629961164
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _27_
timestamp 1629961164
transform -1 0 3772 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629961164
transform -1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_29
timestamp 1629961164
transform 1 0 3772 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_35
timestamp 1629961164
transform 1 0 4324 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _25_
timestamp 1629961164
transform 1 0 4416 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1629961164
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1629961164
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _19_
timestamp 1629961164
transform 1 0 6348 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_66
timestamp 1629961164
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_70
timestamp 1629961164
transform 1 0 7544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_74
timestamp 1629961164
transform 1 0 7912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1629961164
transform -1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1629961164
transform 1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_10
timestamp 1629961164
transform 1 0 2024 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_14
timestamp 1629961164
transform 1 0 2392 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1629961164
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1629961164
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _11_
timestamp 1629961164
transform 1 0 2484 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1629961164
transform -1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1629961164
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_29
timestamp 1629961164
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1629961164
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _26_
timestamp 1629961164
transform -1 0 5796 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_51
timestamp 1629961164
transform 1 0 5796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_55
timestamp 1629961164
transform 1 0 6164 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_57
timestamp 1629961164
transform 1 0 6348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_61
timestamp 1629961164
transform 1 0 6716 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1629961164
transform 1 0 6256 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1629961164
transform -1 0 6716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_74
timestamp 1629961164
transform 1 0 7912 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1629961164
transform -1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _20_
timestamp 1629961164
transform 1 0 7084 0 1 8704
box -38 -48 866 592
<< labels >>
rlabel metal3 s 8935 5720 9735 5840 6 INPUT[0]
port 0 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 INPUT[1]
port 1 nsew signal input
rlabel metal2 s 8298 11079 8354 11879 6 INPUT[2]
port 2 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 INPUT[3]
port 3 nsew signal input
rlabel metal2 s 18 0 74 800 6 INPUT[4]
port 4 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 INPUT[5]
port 5 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 INPUT[6]
port 6 nsew signal input
rlabel metal2 s 5538 11079 5594 11879 6 INPUT[7]
port 7 nsew signal input
rlabel metal3 s 8935 9800 9735 9920 6 INPUT[8]
port 8 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 INPUT[9]
port 9 nsew signal input
rlabel metal2 s 18 11079 74 11879 6 OUTPUT
port 10 nsew signal tristate
rlabel metal5 s 1104 4326 8556 4646 6 VGND
port 11 nsew ground input
rlabel metal5 s 1104 3146 8556 3466 6 VPWR
port 12 nsew power input
rlabel metal2 s 2778 11079 2834 11879 6 clk
port 13 nsew signal input
rlabel metal3 s 8935 1640 9735 1760 6 load
port 14 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 9735 11879
<< end >>
